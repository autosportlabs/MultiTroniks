CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
610 440 30 120 9
20 79 780 560
7 5.000 V
7 5.000 V
3 GND
1000 10
24 100 0 1 0
20 Package,Description,
61 C:\PROGRAM FILES\MICROCODE ENGINEERING\CIRCUITMAKER 6\BOM.DAT
0 7
20 79 780 560
146014226 80
1
37 LVX2 - COMMUNICATION(RS485 & RS422)

49 MULTITRONIKS
1 FREDERICK ROAD
WARREN, NJ. 07059
10 09-17-1998
0
0
60
6 DS8922
94 801 197 0 16 33
0 58 55 19 2 2 2 57 56 43
44 47 48 49 50 46 45
6 DS8922
1 0 2176 0
0
0
0
0
0
0
0
5 DIP16
33

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 1 2 3
4 5 6 7 8 9 10 11 12 13
14 15 16 0
0 0 0 0 1 0 0 0
1 U
8953 0 0
0
0
6 SP232A
94 553 184 0 16 33
0 63 20 62 61 60 59 51 52 57
56 58 55 54 53 2 19
6 SP232A
2 0 4224 0
0
0
0
0
0
0
0
5 DIP16
33

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 1 2 3
4 5 6 7 8 9 10 11 12 13
14 15 16 0
0 0 0 0 1 0 0 0
1 U
4441 0 0
0
0
10 Polar Cap~
219 478 148 0 2 5
0 63 62
0
0 0 320 180
5 0.1uF
-72 -5 -37 3
3 C21
-65 -15 -44 -7
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3618 0 0
0
0
10 Polar Cap~
219 477 178 0 2 5
0 61 60
0
0 0 320 180
5 0.1uF
-70 -3 -35 5
3 C20
-63 -13 -42 -5
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
6153 0 0
0
0
10 Polar Cap~
219 479 100 0 2 5
0 20 19
0
0 0 320 0
5 0.1uF
-65 -7 -30 1
3 C19
-58 -17 -37 -9
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
5394 0 0
0
0
10 Polar Cap~
219 459 234 0 2 5
0 2 59
0
0 0 320 90
5 0.1uF
-53 -6 -18 2
3 C18
-46 -16 -25 -8
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7734 0 0
0
0
7 Ground~
168 459 268 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9914 0 0
0
0
7 Ground~
168 737 259 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3747 0 0
0
0
7 Ground~
168 892 302 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3549 0 0
0
0
10 Polar Cap~
219 650 119 0 2 5
0 19 2
0
0 0 320 270
5 220uF
-16 -34 19 -26
3 C17
-9 -44 12 -36
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7931 0 0
0
0
7 Ground~
168 649 138 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9325 0 0
0
0
10 Capacitor~
219 608 232 0 2 5
0 2 19
0
0 0 320 90
6 0.01uF
-47 10 -5 18
3 C16
-37 0 -16 8
0
0
11 %D %1 %2 %V
0
0
6 CAP0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
8903 0 0
0
0
7 Ground~
168 608 266 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3834 0 0
0
0
6 DS8922
94 795 471 0 16 33
0 36 33 19 2 2 2 35 34 21
23 25 26 27 28 24 22
6 DS8922
3 0 2176 0
0
0
0
0
0
0
0
5 DIP16
33

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 1 2 3
4 5 6 7 8 9 10 11 12 13
14 15 16 0
0 0 0 0 1 0 0 0
1 U
3363 0 0
0
0
6 SP232A
94 554 458 0 16 33
0 42 38 41 40 39 37 29 30 35
34 36 33 32 31 2 19
6 SP232A
4 0 4224 0
0
0
0
0
0
0
0
5 DIP16
33

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 1 2 3
4 5 6 7 8 9 10 11 12 13
14 15 16 0
0 0 0 0 1 0 0 0
1 U
7668 0 0
0
0
10 Polar Cap~
219 476 422 0 2 5
0 42 41
0
0 0 320 180
5 0.1uF
-79 -5 -44 3
3 C15
-72 -15 -51 -7
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
4718 0 0
0
0
10 Polar Cap~
219 474 452 0 2 5
0 40 39
0
0 0 320 180
5 0.1uF
-79 -2 -44 6
3 C14
-72 -12 -51 -4
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3874 0 0
0
0
10 Polar Cap~
219 452 509 0 2 5
0 2 37
0
0 0 320 90
5 0.1uF
-56 -5 -21 3
3 C13
-49 -15 -28 -7
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
6671 0 0
0
0
7 Ground~
168 452 535 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3789 0 0
0
0
7 Ground~
168 741 555 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4871 0 0
0
0
7 Ground~
168 881 571 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3750 0 0
0
0
10 Capacitor~
219 609 515 0 2 5
0 2 19
0
0 0 320 90
6 0.01uF
-49 5 -7 13
3 C12
-39 -5 -18 3
0
0
11 %D %1 %2 %V
0
0
6 CAP0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
8778 0 0
0
0
7 Ground~
168 609 543 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
538 0 0
0
0
10 Capacitor~
219 707 249 0 2 5
0 2 19
0
0 0 320 90
6 0.01uF
-55 -2 -13 6
3 C11
-45 -12 -24 -4
0
0
11 %D %1 %2 %V
0
0
6 CAP0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
6843 0 0
0
0
7 Ground~
168 707 297 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3136 0 0
0
0
10 Polar Cap~
219 491 399 0 2 5
0 38 19
0
0 0 320 0
5 0.1uF
2 -13 37 -5
2 C4
12 -23 26 -15
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
5950 0 0
0
0
10 Capacitor~
219 709 517 0 2 5
0 2 19
0
0 0 320 90
6 0.01uF
-60 -3 -18 5
2 C2
-46 -13 -32 -5
0
0
11 %D %1 %2 %V
0
0
6 CAP0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
5670 0 0
0
0
7 Ground~
168 709 557 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6828 0 0
0
0
7 Ground~
168 64 231 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6735 0 0
0
0
3 DIO
94 427 764 0 2 5
0 7 6
3 DIO
5 0 0 180
12 SINGLE DIODE
-42 -18 42 -10
0
0
0
0
0
0
6 SOT-23
5

0 3 1 3 1 0
0 0 0 0 1 0 0 0
1 D
8365 0 0
0
0
10 SN75ALS180
94 579 652 0 14 29
0 64 65 12 12 6 2 2 66 5
10 67 5 8 8
10 SN75ALS180
6 0 2176 0
0
0
0
0
0
0
0
5 DIP14
29

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 1 2 3 4 5
6 7 8 9 10 11 12 13 14 0
0 0 0 512 1 0 0 0
1 U
4132 0 0
0
0
10 555 Timer~
219 429 728 0 8 17
0 2 6 12 8 11 7 7 8
0
0 0 4416 0
3 555
-11 -36 10 -28
3 X22
-11 -46 10 -38
0
0
29 %D %1 %2 %3 %4 %5 %6 %7 %8 %S
0
0
4 CAN8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
88 0 0 0 1 0 0 0
1 U
4551 0 0
0
0
6 SP232A
94 273 672 0 16 33
0 18 14 17 16 15 13 68 4 6
2 9 69 70 3 2 8
6 SP232A
7 0 6272 0
0
0
0
0
0
0
0
5 DIP16
33

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 1 2 3
4 5 6 7 8 9 10 11 12 13
14 15 16 0
0 0 0 512 1 1 0 0
1 U
3635 0 0
0
0
10 Polar Cap~
219 196 636 0 2 5
0 18 17
0
0 0 320 180
5 0.1uF
-71 -1 -36 7
3 C10
-64 -11 -43 -3
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3973 0 0
0
0
10 Polar Cap~
219 194 666 0 2 5
0 16 15
0
0 0 320 180
5 0.1uF
-70 0 -35 8
2 C9
-60 -10 -46 -2
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3851 0 0
0
0
10 Polar Cap~
219 178 725 0 2 5
0 2 13
0
0 0 320 90
5 0.1uF
-52 -3 -17 5
2 C8
-42 -13 -28 -5
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
8383 0 0
0
0
7 Ground~
168 178 750 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9334 0 0
0
0
10 Capacitor~
219 326 725 0 2 5
0 2 8
0
0 0 320 90
6 0.01uF
-55 6 -13 14
2 C7
-41 -4 -27 4
0
0
11 %D %1 %2 %V
0
0
6 CAP0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7471 0 0
0
0
7 Ground~
168 326 767 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3334 0 0
0
0
7 Ground~
168 516 721 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3559 0 0
0
0
10 Capacitor~
219 555 747 0 2 5
0 2 11
0
0 0 320 180
6 0.01uF
-20 -18 22 -10
2 C6
-6 -28 8 -20
0
0
11 %D %1 %2 %V
0
0
6 CAP0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
984 0 0
0
0
10 Capacitor~
219 513 764 0 2 5
0 2 7
0
0 0 320 180
5 0.1uF
-17 13 18 21
2 C5
-7 3 7 11
0
0
11 %D %1 %2 %V
0
0
6 CAP0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7557 0 0
0
0
7 Ground~
168 610 771 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3146 0 0
0
0
10 Polar Cap~
219 219 609 0 2 5
0 14 8
0
0 0 320 0
5 0.1uF
-93 -6 -58 2
2 C3
-83 -16 -69 -8
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
5687 0 0
0
0
10 Capacitor~
219 628 695 0 2 5
0 2 8
0
0 0 320 90
6 0.01uF
4 -15 46 -7
2 C1
18 -25 32 -17
0
0
11 %D %1 %2 %V
0
0
6 CAP0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7939 0 0
0
0
7 Ground~
168 628 727 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3308 0 0
0
0
6 CON-64
94 137 307 0 64 129
0 2 19 71 72 73 74 75 76 77
78 79 80 81 82 83 84 85 86 87
88 89 90 91 92 3 4 93 94 95
5 10 96 97 98 99 31 32 30 29
100 101 22 24 28 27 26 25 23 21
102 53 54 52 51 103 104 43 44 47
48 49 50 46 45
6 CON-64
8 0 4736 0
0
2 J2
0 -163 14 -155
0
0
0
0
0
0
129

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 21 22 23 24 25 26 27 28 29
30 31 32 33 34 35 36 37 38 39
40 41 42 43 44 45 46 47 48 49
50 51 52 53 54 55 56 57 58 59
60 61 62 63 64 1 2 3 4 5
6 7 8 9 10 11 12 13 14 15
16 17 18 19 20 21 22 23 24 25
26 27 28 29 30 31 32 33 34 35
36 37 38 39 40 41 42 43 44 45
46 47 48 49 50 51 52 53 54 55
56 57 58 59 60 61 62 63 64 0
0 0 0 512 1 0 0 0
1 J
3408 0 0
0
0
9 Resistor~
219 870 137 0 2 5
0 45 19
0
0 0 352 90
2 1k
-18 -6 -4 2
3 R35
-21 -16 0 -8
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9773 0 0
0
0
9 Resistor~
219 895 139 0 2 5
0 43 19
0
0 0 352 90
2 1k
8 -5 22 3
3 R34
5 -15 26 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
691 0 0
0
0
9 Resistor~
219 869 256 0 3 5
0 2 44 -1
0
0 0 352 90
2 1k
8 -5 22 3
3 R33
5 -15 26 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7834 0 0
0
0
9 Resistor~
219 914 257 0 3 5
0 2 46 -1
0
0 0 352 90
2 1k
8 -5 22 3
3 R32
5 -15 26 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3588 0 0
0
0
9 Resistor~
219 865 407 0 2 5
0 22 19
0
0 0 352 90
2 1k
-21 -5 -7 3
3 R31
-24 -15 -3 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4528 0 0
0
0
9 Resistor~
219 884 406 0 2 5
0 21 19
0
0 0 352 90
2 1k
8 -5 22 3
3 R30
5 -15 26 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3303 0 0
0
0
9 Resistor~
219 863 528 0 3 5
0 2 23 -1
0
0 0 352 90
2 1k
8 -5 22 3
3 R29
5 -15 26 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9654 0 0
0
0
9 Resistor~
219 908 524 0 3 5
0 2 24 -1
0
0 0 352 90
2 1k
8 -5 22 3
3 R28
5 -15 26 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9791 0 0
0
0
9 Resistor~
219 360 643 0 2 5
0 9 8
0
0 0 352 90
3 4k7
3 -15 24 -7
3 R27
3 -25 24 -17
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4589 0 0
0
0
9 Resistor~
219 516 689 0 3 5
0 2 12 -1
0
0 0 352 90
3 10k
-19 -9 2 -1
3 R26
-19 -19 2 -11
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
964 0 0
0
0
9 Resistor~
219 488 697 0 2 5
0 8 7
0
0 0 352 270
3 10k
1 -3 22 5
3 R25
1 -13 22 -5
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9151 0 0
0
0
9 Resistor~
219 685 709 0 3 5
0 2 10 -1
0
0 0 352 90
3 4k7
5 -5 26 3
3 R24
5 -15 26 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4745 0 0
0
0
9 Resistor~
219 657 609 0 2 5
0 5 8
0
0 0 352 180
3 4k7
-10 -14 11 -6
3 R23
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8433 0 0
0
0
134
14 25 3 0 0 16512 0 33 47 0 0 6
314 656
349 656
349 784
59 784
59 388
111 388
8 26 4 0 0 8320 0 33 47 0 0 4
232 706
70 706
70 397
111 397
0 30 5 0 0 8320 0 0 47 14 0 5
697 609
697 591
82 591
82 433
111 433
1 0 2 0 0 4096 0 32 0 0 39 2
397 719
338 719
2 0 6 0 0 4096 0 32 0 0 30 2
397 728
379 728
0 1 2 0 0 0 0 0 57 33 0 3
531 679
531 707
516 707
6 0 7 0 0 4096 0 32 0 0 8 2
461 737
488 737
0 0 7 0 0 4096 0 0 0 9 21 2
488 728
488 764
7 2 7 0 0 0 0 32 58 0 0 3
461 728
488 728
488 715
4 0 8 0 0 8192 0 32 0 0 38 3
397 746
390 746
390 609
1 1 2 0 0 0 0 45 46 0 0 2
628 704
628 721
0 2 8 0 0 0 0 0 45 38 0 2
628 634
628 686
11 1 9 0 0 4224 0 33 56 0 0 3
314 686
360 686
360 661
0 1 5 0 0 0 0 0 60 16 0 4
650 643
697 643
697 609
675 609
0 2 8 0 0 0 0 0 60 38 0 2
627 609
639 609
9 12 5 0 0 0 0 31 31 0 0 4
611 670
650 670
650 643
611 643
14 0 8 0 0 0 0 31 0 0 38 2
611 625
628 625
0 2 10 0 0 4096 0 0 59 19 0 2
685 661
685 691
10 31 10 0 0 12416 0 31 47 0 0 6
611 661
685 661
685 579
95 579
95 442
111 442
0 1 2 0 0 4096 0 0 59 24 0 3
610 764
685 764
685 727
2 1 7 0 0 4224 0 42 30 0 0 2
504 764
435 764
2 5 11 0 0 4224 0 41 32 0 0 3
546 747
461 747
461 746
1 0 2 0 0 0 0 41 0 0 24 3
564 747
610 747
610 755
1 1 2 0 0 4096 0 42 43 0 0 5
522 764
610 764
610 755
610 755
610 765
1 0 8 0 0 0 0 58 0 0 32 3
488 679
488 672
471 672
1 1 2 0 0 0 0 57 40 0 0 2
516 707
516 715
2 0 12 0 0 4096 0 57 0 0 28 2
516 671
516 652
4 0 12 0 0 4096 0 31 0 0 29 3
547 652
516 652
516 643
3 3 12 0 0 4224 0 31 32 0 0 4
547 643
370 643
370 737
397 737
0 2 6 0 0 4096 0 0 30 35 0 3
379 706
379 764
412 764
10 0 2 0 0 0 0 33 0 0 39 2
314 696
338 696
8 0 8 0 0 0 0 32 0 0 38 3
461 719
471 719
471 609
7 6 2 0 0 0 0 31 31 0 0 4
547 679
530 679
530 670
547 670
2 0 8 0 0 0 0 56 0 0 38 2
360 625
360 609
9 5 6 0 0 12416 0 33 31 0 0 4
314 706
379 706
379 661
547 661
0 2 8 0 0 0 0 0 38 37 0 2
326 636
326 716
16 0 8 0 0 0 0 33 0 0 38 3
314 636
326 636
326 609
2 13 8 0 0 4224 0 44 31 0 0 4
225 609
628 609
628 634
611 634
0 15 2 0 0 8192 0 0 33 40 0 4
326 736
338 736
338 646
314 646
1 1 2 0 0 0 0 39 38 0 0 2
326 761
326 734
1 1 2 0 0 0 0 37 36 0 0 2
178 744
178 734
2 6 13 0 0 8320 0 36 33 0 0 3
178 717
178 686
232 686
2 1 14 0 0 4224 0 33 44 0 0 4
232 646
177 646
177 609
208 609
2 5 15 0 0 12416 0 35 33 0 0 4
184 666
160 666
160 676
232 676
4 1 16 0 0 4224 0 33 35 0 0 2
232 666
201 666
2 3 17 0 0 12416 0 34 33 0 0 4
186 636
160 636
160 656
232 656
1 1 18 0 0 4224 0 33 34 0 0 2
232 636
203 636
1 1 2 0 0 0 0 29 47 0 0 3
64 225
64 172
111 172
2 0 19 0 0 4096 0 27 0 0 97 2
709 508
709 456
1 1 2 0 0 0 0 28 27 0 0 2
709 551
709 526
15 0 2 0 0 8320 0 15 0 0 57 4
595 432
625 432
625 531
609 531
2 0 19 0 0 4096 0 22 0 0 97 2
609 506
609 422
0 0 19 0 0 0 0 0 0 134 118 2
626 148
626 100
2 0 19 0 0 0 0 12 0 0 134 2
608 223
608 148
0 2 19 0 0 8320 0 0 47 118 0 5
564 100
564 81
85 81
85 181
111 181
1 2 20 0 0 12416 0 5 2 0 0 4
468 100
453 100
453 158
512 158
1 1 2 0 0 0 0 22 23 0 0 2
609 524
609 537
9 1 21 0 0 8192 0 14 53 0 0 3
827 501
884 501
884 424
0 1 22 0 0 8192 0 0 52 67 0 3
866 438
865 438
865 425
6 0 2 0 0 0 0 14 0 0 84 2
763 483
741 483
15 0 2 0 0 0 0 2 0 0 110 4
594 158
626 158
626 251
608 251
2 0 19 0 0 0 0 24 0 0 134 2
707 240
707 182
1 1 2 0 0 0 0 25 24 0 0 2
707 291
707 258
0 0 19 0 0 0 0 0 0 118 80 2
694 100
694 382
0 49 21 0 0 16512 0 0 47 58 0 5
884 501
884 500
977 500
977 307
177 307
0 48 23 0 0 12416 0 0 47 78 0 4
862 492
969 492
969 316
177 316
16 42 22 0 0 12416 0 14 47 0 0 4
827 438
914 438
914 370
177 370
0 43 24 0 0 12416 0 0 47 77 0 4
908 447
924 447
924 361
177 361
11 47 25 0 0 12416 0 14 47 0 0 4
827 483
961 483
961 325
177 325
12 46 26 0 0 12416 0 14 47 0 0 4
827 474
952 474
952 334
177 334
13 45 27 0 0 12416 0 14 47 0 0 4
827 465
942 465
942 343
177 343
14 44 28 0 0 12416 0 14 47 0 0 4
827 456
933 456
933 352
177 352
7 39 29 0 0 4224 0 15 47 0 0 4
513 482
278 482
278 397
177 397
8 38 30 0 0 4224 0 15 47 0 0 4
513 492
268 492
268 406
177 406
14 36 31 0 0 12416 0 15 47 0 0 6
595 442
647 442
647 565
245 565
245 424
177 424
13 37 32 0 0 12416 0 15 47 0 0 6
595 452
637 452
637 556
256 556
256 415
177 415
15 2 24 0 0 0 0 14 55 0 0 3
827 447
908 447
908 506
10 2 23 0 0 0 0 14 54 0 0 3
827 492
863 492
863 510
2 0 19 0 0 0 0 52 0 0 80 2
865 389
865 382
2 0 19 0 0 0 0 53 0 0 91 4
884 388
884 382
694 382
694 400
1 0 2 0 0 0 0 21 0 0 82 2
881 565
881 553
1 1 2 0 0 0 0 54 55 0 0 4
863 546
863 553
908 553
908 542
5 0 2 0 0 0 0 14 0 0 84 2
763 474
741 474
1 4 2 0 0 0 0 20 14 0 0 3
741 549
741 465
763 465
12 2 33 0 0 4224 0 15 14 0 0 4
595 462
684 462
684 447
763 447
10 8 34 0 0 4224 0 15 14 0 0 4
595 482
725 482
725 501
763 501
9 7 35 0 0 4224 0 15 14 0 0 2
595 492
763 492
11 1 36 0 0 4224 0 15 14 0 0 4
595 472
724 472
724 438
763 438
1 1 2 0 0 0 0 19 18 0 0 2
452 529
452 518
2 6 37 0 0 8320 0 18 15 0 0 3
452 501
452 472
513 472
2 0 19 0 0 0 0 26 0 0 97 4
497 399
497 400
694 400
694 422
2 1 38 0 0 4224 0 15 26 0 0 4
513 432
452 432
452 399
480 399
2 5 39 0 0 12416 0 17 15 0 0 4
464 452
437 452
437 462
513 462
4 1 40 0 0 4224 0 15 17 0 0 2
513 452
481 452
2 3 41 0 0 12416 0 16 15 0 0 4
466 422
444 422
444 442
513 442
1 1 42 0 0 4224 0 15 16 0 0 2
513 422
483 422
16 3 19 0 0 0 0 15 14 0 0 4
595 422
694 422
694 456
763 456
0 57 43 0 0 12416 0 0 47 115 0 6
895 227
983 227
983 18
255 18
255 235
177 235
0 58 44 0 0 12416 0 0 47 114 0 6
868 218
975 218
975 26
245 26
245 226
177 226
0 64 45 0 0 12416 0 0 47 116 0 6
870 164
920 164
920 72
190 72
190 172
177 172
0 63 46 0 0 12416 0 0 47 113 0 6
914 173
930 173
930 64
199 64
199 181
177 181
11 59 47 0 0 12416 0 1 47 0 0 6
833 209
967 209
967 34
237 34
237 217
177 217
12 60 48 0 0 12416 0 1 47 0 0 6
833 200
958 200
958 42
226 42
226 208
177 208
13 61 49 0 0 12416 0 1 47 0 0 6
833 191
948 191
948 49
218 49
218 199
177 199
14 62 50 0 0 12416 0 1 47 0 0 6
833 182
939 182
939 57
208 57
208 190
177 190
7 54 51 0 0 4224 0 2 47 0 0 4
512 208
270 208
270 262
177 262
8 53 52 0 0 4224 0 2 47 0 0 4
512 218
279 218
279 271
177 271
14 51 53 0 0 12416 0 2 47 0 0 4
594 168
645 168
645 289
177 289
13 52 54 0 0 12416 0 2 47 0 0 4
594 178
637 178
637 280
177 280
1 1 2 0 0 0 0 13 12 0 0 2
608 260
608 241
1 2 2 0 0 0 0 11 10 0 0 4
649 132
649 122
649 122
649 126
1 0 19 0 0 0 0 10 0 0 118 2
649 109
649 100
15 2 46 0 0 0 0 1 51 0 0 3
833 173
914 173
914 239
10 2 44 0 0 0 0 1 50 0 0 3
833 218
869 218
869 238
9 1 43 0 0 0 0 1 49 0 0 3
833 227
895 227
895 157
16 1 45 0 0 0 0 1 48 0 0 3
833 164
870 164
870 155
2 0 19 0 0 0 0 48 0 0 118 3
870 119
871 119
871 100
2 2 19 0 0 0 0 49 5 0 0 3
895 121
895 100
485 100
1 0 2 0 0 0 0 9 0 0 120 2
892 296
892 286
1 1 2 0 0 0 0 50 51 0 0 4
869 274
869 286
914 286
914 275
6 0 2 0 0 0 0 1 0 0 123 2
769 209
737 209
5 0 2 0 0 0 0 1 0 0 123 2
769 200
737 200
1 4 2 0 0 0 0 8 1 0 0 3
737 253
737 191
769 191
12 2 55 0 0 12416 0 2 1 0 0 4
594 188
655 188
655 173
769 173
10 8 56 0 0 4224 0 2 1 0 0 4
594 208
719 208
719 227
769 227
9 7 57 0 0 4224 0 2 1 0 0 2
594 218
769 218
11 1 58 0 0 4224 0 2 1 0 0 4
594 198
720 198
720 164
769 164
1 1 2 0 0 0 0 7 6 0 0 2
459 262
459 243
2 6 59 0 0 8320 0 6 2 0 0 3
459 226
459 198
512 198
2 5 60 0 0 12416 0 4 2 0 0 4
467 178
443 178
443 188
512 188
4 1 61 0 0 4224 0 2 4 0 0 2
512 178
484 178
2 3 62 0 0 12416 0 3 2 0 0 4
468 148
443 148
443 168
512 168
1 1 63 0 0 4224 0 2 3 0 0 2
512 148
485 148
16 3 19 0 0 0 0 2 1 0 0 4
594 148
665 148
665 182
769 182
12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
107 561 123 585
111 565 119 581
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
89 587 105 611
93 591 101 607
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
70 372 94 396
74 376 90 392
2 RD
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
75 394 99 418
79 398 95 414
2 TD
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
277 559 309 583
281 563 305 579
3 RTS
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
265 539 297 563
269 543 293 559
3 CTS
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
216 384 240 408
220 388 236 404
2 RD
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
269 484 293 508
273 488 289 504
2 TD
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
330 284 362 308
334 288 358 304
3 RTS
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
299 266 331 290
303 270 327 286
3 CTS
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
279 212 303 236
283 216 299 232
2 TD
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
213 247 237 271
217 251 233 267
2 RD
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
