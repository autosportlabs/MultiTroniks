CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 10 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 190 30 100 9
21 78 780 559
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 1 1 0
20 Package,Description,
61 C:\PROGRAM FILES\MICROCODE ENGINEERING\CIRCUITMAKER 6\BOM.DAT
0 7
21 78 780 559
146276370 80
2
41 Title:3 PHASE /208Y/120VAC WIRING DIAGRAM
51 MULTITRONIKS
ONE FREDERICK ROAD, WARREN, NJ 07059.
8 02-22-99
0
4 LVX2
49
5 Ter1~
94 246 271 0 1 3
0 40
5 Ter1~
1 0 0 180
0
3 U39
-10 -16 11 -8
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 J
8953 0 0
0
0
5 Ter1~
94 246 281 0 1 3
0 38
5 Ter1~
2 0 0 180
0
3 U38
-10 -16 11 -8
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 J
4441 0 0
0
0
5 Ter1~
94 245 325 0 1 3
0 7
5 Ter1~
3 0 0 180
0
3 U37
-10 -16 11 -8
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 J
3618 0 0
0
0
5 Ter1~
94 245 335 0 1 3
0 6
5 Ter1~
4 0 0 180
0
3 U36
2 -17 23 -9
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 J
6153 0 0
0
0
5 Ter1~
94 245 345 0 1 3
0 5
5 Ter1~
5 0 0 180
0
3 U35
-12 -15 9 -7
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 J
5394 0 0
0
0
5 Ter1~
94 245 355 0 1 3
0 36
5 Ter1~
6 0 0 180
0
3 U34
-10 -16 11 -8
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 J
7734 0 0
0
0
5 Ter1~
94 404 334 0 1 3
0 40
5 Ter1~
7 0 0 270
0
3 U33
-12 -23 9 -15
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 J
9914 0 0
0
0
5 Ter1~
94 423 334 0 1 3
0 39
5 Ter1~
8 0 0 270
0
3 U32
-12 -23 9 -15
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 J
3747 0 0
0
0
5 Ter1~
94 443 335 0 1 3
0 38
5 Ter1~
9 0 0 270
0
3 U31
-12 -23 9 -15
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 J
3549 0 0
0
0
5 Ter1~
94 404 252 0 1 3
0 42
5 Ter1~
10 0 0 90
0
3 U30
8 -3 29 5
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 J
7931 0 0
0
0
5 Ter1~
94 423 252 0 1 3
0 43
5 Ter1~
11 0 0 90
0
3 U29
8 -3 29 5
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 J
9325 0 0
0
0
5 Ter1~
94 441 252 0 1 3
0 44
5 Ter1~
12 0 0 90
0
3 U28
8 -3 29 5
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 J
8903 0 0
0
0
5 Ter1~
94 553 610 0 1 3
0 54
5 Ter1~
13 0 0 270
0
3 U27
-12 -23 9 -15
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 J
3834 0 0
0
0
5 Ter1~
94 574 610 0 1 3
0 55
5 Ter1~
14 0 0 270
0
3 U26
-12 -23 9 -15
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 J
3363 0 0
0
0
5 Ter1~
94 597 610 0 1 3
0 56
5 Ter1~
15 0 0 270
0
3 U25
-12 -23 9 -15
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 J
7668 0 0
0
0
5 Ter1~
94 553 512 0 1 3
0 45
5 Ter1~
16 0 0 90
0
3 U24
8 -3 29 5
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 J
4718 0 0
0
0
5 Ter1~
94 578 513 0 1 3
0 46
5 Ter1~
17 0 0 90
0
3 U23
8 -3 29 5
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 J
3874 0 0
0
0
5 Ter1~
94 603 512 0 1 3
0 31
5 Ter1~
18 0 0 90
0
3 U22
8 -3 29 5
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 J
6671 0 0
0
0
5 Ter1~
94 683 121 0 1 3
0 44
5 Ter1~
19 0 0 602
0
3 U21
8 -3 29 5
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 J
3789 0 0
0
0
5 Ter1~
94 656 121 0 1 3
0 43
5 Ter1~
20 0 0 602
0
3 U20
8 -3 29 5
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 J
4871 0 0
0
0
5 Ter1~
94 628 121 0 1 3
0 42
5 Ter1~
21 0 0 602
0
3 U19
8 -3 29 5
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 J
3750 0 0
0
0
5 Ter1~
94 690 224 0 1 3
0 59
5 Ter1~
22 0 0 782
0
3 U18
-12 -23 9 -15
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 J
8778 0 0
0
0
5 Ter1~
94 674 224 0 1 3
0 35
5 Ter1~
23 0 0 782
0
3 U17
-12 -23 9 -15
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 J
538 0 0
0
0
5 Ter1~
94 659 224 0 1 3
0 29
5 Ter1~
24 0 0 782
0
3 U16
-12 -23 9 -15
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 J
6843 0 0
0
0
5 Ter1~
94 642 224 0 1 3
0 26
5 Ter1~
25 0 0 782
0
3 U15
-12 -23 9 -15
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 J
3136 0 0
0
0
5 Ter1~
94 626 224 0 1 3
0 60
5 Ter1~
26 0 0 782
0
3 U14
-12 -23 9 -15
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 J
5950 0 0
0
0
10 TER BLOCK~
94 554 390 0 2 5
0 45 29
10 TER BLOCK~
27 0 0 90
0
3 U13
7 -7 28 1
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 0 1 0 0 0
1 J
5670 0 0
0
0
10 TER BLOCK~
94 719 394 0 2 5
0 36 8
10 TER BLOCK~
28 0 0 90
0
3 U11
7 -7 28 1
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 0 1 0 0 0
1 J
6828 0 0
0
0
10 TER BLOCK~
94 709 394 0 2 5
0 37 26
10 TER BLOCK~
29 0 0 90
0
3 U10
7 -7 28 1
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 0 1 0 0 0
1 J
6735 0 0
0
0
10 TER BLOCK~
94 579 391 0 2 5
0 46 35
10 TER BLOCK~
30 0 0 90
0
2 U9
8 -7 22 1
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 0 1 0 0 0
1 J
8365 0 0
0
0
10 TER BLOCK~
94 589 391 0 2 5
0 34 63
10 TER BLOCK~
31 0 0 90
0
2 U8
8 -7 22 1
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
1 J
4132 0 0
0
0
10 TER BLOCK~
94 607 392 0 2 5
0 31 59
10 TER BLOCK~
32 0 0 90
0
2 U6
8 -7 22 1
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 0 1 0 0 0
1 J
4551 0 0
0
0
10 TER BLOCK~
94 626 392 0 2 5
0 9 60
10 TER BLOCK~
33 0 0 90
0
2 U5
8 -7 22 1
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 0 1 0 0 0
1 J
3635 0 0
0
0
10 TER BLOCK~
94 636 392 0 2 5
0 33 64
10 TER BLOCK~
34 0 0 90
0
2 U4
8 -7 22 1
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
1 J
3973 0 0
0
0
10 TER BLOCK~
94 655 393 0 2 5
0 56 10
10 TER BLOCK~
35 0 0 90
0
2 U3
8 -7 22 1
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 0 1 0 0 0
1 J
3851 0 0
0
0
10 TER BLOCK~
94 673 393 0 2 5
0 55 11
10 TER BLOCK~
36 0 0 90
0
2 U2
8 -7 22 1
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 0 1 0 0 0
1 J
8383 0 0
0
0
10 TER BLOCK~
94 691 394 0 2 5
0 54 12
10 TER BLOCK~
37 0 0 90
0
2 U1
8 -7 22 1
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 0 1 0 0 0
1 J
9334 0 0
0
0
5 Ter1~
94 81 325 0 1 3
0 2
5 Ter1~
38 0 0 270
0
3 U42
-12 -23 9 -15
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 J
7471 0 0
0
0
5 Ter1~
94 91 325 0 1 3
0 3
5 Ter1~
39 0 0 270
0
3 U41
-12 -23 9 -15
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 J
3334 0 0
0
0
5 Ter1~
94 101 325 0 1 3
0 4
5 Ter1~
40 0 0 270
0
3 U40
-12 -23 9 -15
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 J
3559 0 0
0
0
5 Ter1~
94 86 373 0 1 3
0 38
5 Ter1~
41 0 0 270
0
3 U45
-12 -23 9 -15
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 J
984 0 0
0
0
5 Ter1~
94 76 373 0 1 3
0 39
5 Ter1~
42 0 0 270
0
3 U46
-12 -23 9 -15
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 J
7557 0 0
0
0
5 Ter1~
94 67 373 0 1 3
0 40
5 Ter1~
43 0 0 270
0
3 U47
-12 -23 9 -15
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 J
3146 0 0
0
0
5 Ter1~
94 58 325 0 1 3
0 38
5 Ter1~
44 0 0 270
0
3 U48
-12 -23 9 -15
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 J
5687 0 0
0
0
5 Ter1~
94 48 325 0 1 3
0 40
5 Ter1~
45 0 0 270
0
3 U49
-12 -23 9 -15
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 J
7939 0 0
0
0
5 Ter1~
94 32 353 0 1 3
0 37
5 Ter1~
46 0 0 270
0
3 U50
-12 -23 9 -15
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 J
3308 0 0
0
0
5 Ter1~
94 121 351 0 1 3
0 36
5 Ter1~
47 0 0 270
0
3 U51
-12 -23 9 -15
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 J
3408 0 0
0
0
5 Fuse~
219 904 280 0 2 5
0 34 32
0
0 0 4416 0
3 10A
-7 -19 14 -11
2 F1
-7 -26 7 -18
0
0
11 %D %1 %2 %S
0
23 alias:XFUSE {CURRENT=1}
4 FUSE
5

0 1 2 1 2 0
88 0 0 0 1 0 0 0
1 F
9773 0 0
0
0
7 L21-30P
94 927 398 0 1 3
0 0
7 L21-30P
48 0 0 0
0
2 C2
-3 -58 11 -50
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
1 C
691 0 0
0
0
67
1 0 2 0 0 20608 0 38 0 0 0 6
81 339
81 348
101 348
101 397
147 397
147 159
1 0 3 0 0 20608 0 39 0 0 0 6
91 339
91 344
105 344
105 392
142 392
142 160
1 0 4 0 0 16512 0 40 0 0 0 5
101 339
109 339
109 388
138 388
138 158
1 0 5 0 0 8320 0 5 0 0 0 3
228 346
186 346
186 218
1 0 6 0 0 8320 0 4 0 0 0 3
228 336
192 336
192 217
1 0 7 0 0 8320 0 3 0 0 0 3
228 326
199 326
199 217
2 0 8 0 0 12416 0 28 0 0 0 7
717 376
719 376
719 372
913 372
913 388
929 388
929 398
1 0 9 0 0 8320 0 33 0 0 0 5
624 407
624 446
863 446
863 399
895 399
2 0 10 0 0 8320 0 35 0 0 0 6
653 375
653 332
1007 332
1007 455
930 455
930 434
2 0 11 0 0 8320 0 36 0 0 0 5
671 375
671 339
990 339
990 400
967 400
2 0 12 0 0 8320 0 37 0 0 0 4
689 376
689 347
930 347
930 363
0 0 13 0 0 8320 0 0 0 0 0 3
125 461
125 488
92 488
0 0 14 0 0 4224 0 0 0 0 0 3
255 442
255 505
224 505
0 0 15 0 0 4224 0 0 0 0 0 3
401 403
401 494
379 494
0 0 16 0 0 4224 0 0 0 0 0 3
415 422
415 494
379 494
0 0 17 0 0 4224 0 0 0 0 0 3
2 488
106 488
106 454
0 0 18 0 0 4224 0 0 0 0 0 3
233 415
233 505
152 505
0 0 19 0 0 8320 0 0 0 0 0 3
432 433
432 494
301 494
0 0 20 0 0 12416 0 0 0 0 0 4
474 278
519 278
519 309
607 309
0 0 21 0 0 12416 0 0 0 0 0 4
473 278
525 278
525 301
580 301
0 0 22 0 0 12416 0 0 0 0 0 4
438 177
473 177
473 160
541 160
0 0 23 0 0 12416 0 0 0 0 0 4
418 145
448 145
448 160
501 160
0 0 24 0 0 4224 0 0 0 0 0 2
399 160
484 160
0 0 25 0 0 12416 0 0 0 0 0 4
636 315
717 315
717 302
813 302
0 0 27 0 0 4224 0 0 0 0 0 2
627 256
557 256
0 0 28 0 0 4224 0 0 0 0 0 2
555 278
471 278
1 2 26 0 0 4224 0 25 29 0 0 4
640 238
640 327
707 327
707 376
1 2 29 0 0 8320 0 24 27 0 0 4
657 238
657 274
552 274
552 372
0 0 30 0 0 4224 0 0 0 0 0 3
954 270
1028 270
1028 315
2 0 8 0 0 0 0 28 0 0 0 5
717 376
717 325
862 325
862 313
1022 313
1 1 31 0 0 4224 0 32 18 0 0 4
605 407
605 482
602 482
602 497
2 0 32 0 0 12416 0 48 0 0 0 4
926 280
929 280
929 294
1020 294
1 0 33 0 0 8320 0 34 0 0 0 5
634 407
634 427
851 427
851 304
1021 304
1 1 34 0 0 8320 0 31 48 0 0 5
587 406
587 437
842 437
842 280
882 280
2 1 35 0 0 8320 0 30 23 0 0 4
577 373
577 283
672 283
672 238
1 1 36 0 0 8320 0 28 47 0 0 4
717 409
717 463
121 463
121 365
1 1 37 0 0 8320 0 46 29 0 0 4
32 367
32 454
707 454
707 409
1 1 38 0 0 12416 0 9 44 0 0 5
443 349
447 349
447 444
58 444
58 339
1 1 38 0 0 0 0 9 41 0 0 4
443 349
443 433
86 433
86 387
1 1 39 0 0 8320 0 8 42 0 0 4
423 348
423 424
76 424
76 387
1 1 40 0 0 12416 0 7 45 0 0 5
404 348
409 348
409 415
48 415
48 339
1 1 40 0 0 0 0 7 43 0 0 4
404 348
404 405
67 405
67 387
0 0 41 0 0 12416 0 0 0 0 0 7
26 210
26 192
131 192
131 380
26 380
26 192
28 192
1 1 36 0 0 0 0 6 28 0 0 6
228 356
192 356
192 472
719 472
719 409
717 409
1 1 38 0 0 0 0 9 2 0 0 6
443 349
439 349
439 386
205 386
205 282
229 282
1 1 40 0 0 0 0 7 1 0 0 6
404 348
400 348
400 395
213 395
213 272
229 272
1 1 42 0 0 8320 0 10 21 0 0 4
403 237
403 75
627 75
627 106
1 1 43 0 0 8320 0 20 11 0 0 4
655 106
655 84
422 84
422 237
1 1 44 0 0 8320 0 12 19 0 0 4
440 237
440 93
682 93
682 106
1 1 45 0 0 4224 0 16 27 0 0 2
552 497
552 405
1 1 46 0 0 4224 0 17 30 0 0 2
577 498
577 406
0 0 47 0 0 4224 0 0 0 0 0 2
698 368
698 413
0 0 48 0 0 4224 0 0 0 0 0 2
680 368
680 415
0 0 49 0 0 4224 0 0 0 0 0 2
662 366
662 416
0 0 50 0 0 4224 0 0 0 0 0 2
643 367
643 418
0 0 51 0 0 4224 0 0 0 0 0 2
614 366
614 418
0 0 52 0 0 4224 0 0 0 0 0 2
596 366
596 418
0 0 53 0 0 4224 0 0 0 0 0 2
564 366
564 419
1 1 54 0 0 4224 0 37 13 0 0 4
689 409
689 653
553 653
553 624
1 1 55 0 0 4224 0 36 14 0 0 4
671 408
671 641
574 641
574 624
1 1 56 0 0 4224 0 35 15 0 0 4
653 408
653 630
597 630
597 624
0 0 57 0 0 8320 0 0 0 0 0 6
578 503
616 503
616 617
535 617
535 503
578 503
0 0 58 0 0 12416 0 0 0 0 0 6
389 261
389 243
455 243
455 342
389 342
389 243
2 1 59 0 0 8320 0 32 22 0 0 4
605 374
605 304
688 304
688 238
2 1 60 0 0 4224 0 33 26 0 0 2
624 374
624 238
0 0 61 0 0 12416 0 0 0 0 0 6
700 116
700 231
612 231
612 111
700 111
700 116
0 0 62 0 0 4224 0 0 0 0 0 5
234 157
234 376
348 376
348 157
234 157
49
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 9
716 291 793 312
720 295 790 310
9 GRN 12SWG
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
929 440 953 464
933 444 949 460
2 L3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
975 386 999 410
979 390 995 406
2 L2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
907 340 931 364
911 344 927 360
2 L1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
929 377 945 401
933 381 941 397
1 G
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
868 387 884 411
872 391 880 407
1 N
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
121 124 177 168
125 128 173 160
11 TO Y
MOTOR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
173 181 229 225
177 185 225 217
11 TO X
MOTOR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
787 361 837 382
790 364 832 379
5 GREEN
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
836 436 886 457
840 439 882 454
5 WHITE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
827 461 1018 482
831 464 1014 479
22 4POLE 5-WIRE GROUNDING
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 9
386 283 456 304
390 287 453 302
9 CONTACTOR
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 9
301 484 368 504
304 487 364 501
9 BLK 16SWG
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
51 294 67 315
54 298 62 313
1 t
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
39 294 55 315
43 298 51 313
1 r
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
72 296 88 317
76 299 84 314
1 U
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
83 296 99 317
86 299 94 314
1 V
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
92 296 108 317
96 299 104 314
1 W
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
58 345 74 366
62 348 70 363
1 R
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
68 345 84 366
71 348 79 363
1 S
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
77 344 93 365
81 348 89 363
1 T
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
112 323 128 344
116 326 124 341
1 E
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
24 325 40 346
27 328 35 343
1 E
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
252 345 268 366
255 349 263 364
1 E
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
254 272 270 293
257 275 265 290
1 T
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
253 262 269 283
256 265 264 280
1 R
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
251 335 267 356
255 338 263 353
1 W
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
251 325 267 346
255 328 263 343
1 V
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
253 315 269 336
256 318 264 333
1 U
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 9
946 283 1013 303
949 286 1009 300
9 BLK 16SWG
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 9
946 293 1013 313
949 296 1009 310
9 WHT 16SWG
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 9
945 303 1012 323
948 306 1008 320
9 GRN 16SWG
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 12
950 248 1037 268
954 251 1034 265
12 TO ON/OFF SW
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 9
950 259 1017 279
953 262 1013 276
9 TOP FRAME
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
633 158 680 178
637 162 677 176
6 FILTER
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
617 196 631 216
620 199 627 213
1 N
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
618 127 632 147
622 131 629 145
1 R
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
646 127 660 147
650 130 657 144
1 S
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
674 128 688 148
677 131 684 145
1 T
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
682 196 696 216
685 199 692 213
1 T
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
633 195 647 215
637 199 644 213
1 E
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
665 196 679 216
668 199 675 213
1 S
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
650 196 664 216
654 199 661 213
1 R
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 9
549 240 616 260
553 243 613 257
9 WHT 12SWG
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 9
476 150 543 170
480 153 540 167
9 BLK 12SWG
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 9
469 267 536 287
473 270 533 284
9 BLK 12SWG
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 9
14 478 81 498
18 481 78 495
9 GRN 16SWG
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 10
147 494 221 514
151 497 218 511
10 BRN 16 SWG
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
555 544 595 568
559 548 591 564
4 MCCB
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
