CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
70 20 30 100 9
0 66 1024 740
7 5.000 V
7 5.000 V
3 GND
1000 10
24 100 0 1 0
20 Package,Description,
61 C:\PROGRAM FILES\MICROCODE ENGINEERING\CIRCUITMAKER 6\BOM.DAT
0 7
0 66 1024 740
9961490 0
0
0
0
0
0
0
16
7 Ground~
168 701 570 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8953 0 0
0
0
7 Ground~
168 661 254 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4441 0 0
0
0
7 Ground~
168 670 473 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3618 0 0
0
0
7 Ground~
168 661 124 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6153 0 0
0
0
7 Ground~
168 492 306 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5394 0 0
0
0
7 Ground~
168 221 211 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7734 0 0
0
0
7 Ground~
168 231 472 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9914 0 0
0
0
4 2003
94 448 264 0 16 33
0 15 25 26 27 28 29 14 2 12
30 31 32 33 34 10 11
4 2003
1 0 6528 512
2 U1
-8 -55 6 -47
2 U1
-8 -65 6 -57
0
0
0
0
0
5 DIP16
33

0 1 2 3 4 5 6 7 8 16
15 14 13 12 11 10 9 1 2 3
4 5 6 7 8 16 15 14 13 12
11 10 9 0
0 0 0 512 1 1 0 0
1 A
3747 0 0
0
0
4 CON9
94 194 438 0 9 19
0 20 19 18 17 16 7 2 12 11
4 CON9
2 0 4736 0
2 J2
-31 -100 -17 -92
2 J2
-36 -99 -22 -91
0
0
0
0
0
4 SIP9
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
0 0 0 0 1 0 0 0
1 A
3549 0 0
0
0
5 CON12
94 191 188 0 12 25
0 24 23 22 21 13 8 2 10 11
35 36 37
5 CON12
3 0 4480 0
2 J1
-36 -109 -22 -101
2 J1
-31 -120 -17 -112
0
0
0
0
0
5 SIP12
25

0 1 2 3 4 5 6 7 8 9
10 11 12 1 2 3 4 5 6 7
8 9 10 11 12 0
0 0 0 512 1 0 0 0
1 A
7931 0 0
0
0
5 CON12
94 766 413 0 12 25
0 2 24 23 22 21 2 2 20 19
18 17 2
5 CON12
4 0 4480 512
2 J5
-25 -110 -11 -102
2 J5
-31 -120 -17 -112
0
0
0
0
0
5 SIP12
25

0 1 2 3 4 5 6 7 8 9
10 11 12 1 2 3 4 5 6 7
8 9 10 11 12 0
0 0 0 0 1 0 0 0
1 A
9325 0 0
0
0
4 CON2
94 708 109 0 2 5
0 11 9
4 CON2
5 0 4480 512
2 J3
-6 -29 8 -21
2 J3
-11 -40 3 -32
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 A
8903 0 0
0
0
5 CON10
94 715 236 0 10 21
0 13 14 16 15 38 2 8 2 7
39
5 CON10
6 0 4480 0
2 J4
-17 -60 -3 -52
2 J4
-17 -70 -3 -62
0
0
0
0
0
5 IDC10
21

0 2 4 6 8 10 1 3 5 7
9 2 4 6 8 10 1 3 5 7
9 0
0 0 0 512 1 0 0 0
1 A
3834 0 0
0
0
4 CON5
94 746 527 0 5 11
0 3 4 5 6 2
4 CON5
7 0 4480 0
2 J8
-7 -42 7 -34
0
0
0
0
0
0
0
11

0 1 2 3 4 5 1 2 3 4
5 0
0 0 0 0 1 0 0 0
1 J
3363 0 0
0
0
4 CON2
94 180 516 0 2 5
0 3 4
4 CON2
8 0 4480 0
2 J6
-16 -30 -2 -22
0
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 A
7668 0 0
0
0
4 CON2
94 182 600 0 2 5
0 5 6
4 CON2
9 0 4480 0
2 J7
-16 -30 -2 -22
0
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 A
4718 0 0
0
0
35
1 1 3 0 0 4224 0 15 14 0 0 2
187 506
724 506
2 2 4 0 0 4224 0 14 15 0 0 2
724 516
187 516
1 3 5 0 0 12416 0 16 14 0 0 4
189 590
293 590
293 526
724 526
4 2 6 0 0 4224 0 14 16 0 0 4
724 536
303 536
303 600
189 600
1 5 2 0 0 8192 0 1 14 0 0 3
701 564
701 546
724 546
8 0 2 0 0 0 0 13 0 0 7 2
673 217
661 217
6 1 2 0 0 8192 0 13 2 0 0 3
673 196
661 196
661 248
6 9 7 0 0 12416 0 9 13 0 0 6
187 408
228 408
228 319
575 319
575 226
673 226
6 7 8 0 0 12416 0 10 13 0 0 4
184 148
416 148
416 206
673 206
0 2 9 0 0 4224 0 0 12 0 0 3
688 110
688 109
687 109
8 15 10 0 0 12416 0 10 8 0 0 4
184 168
259 168
259 288
415 288
0 1 2 0 0 0 0 0 4 0 0 3
685 109
661 109
661 118
0 9 11 0 0 8192 0 0 9 14 0 4
391 298
191 298
191 438
187 438
0 16 11 0 0 0 0 0 8 15 0 3
391 178
391 298
415 298
1 9 11 0 0 4224 0 12 10 0 0 4
687 99
391 99
391 178
184 178
8 9 12 0 0 12416 0 9 8 0 0 4
187 428
202 428
202 228
415 228
1 5 13 0 0 12416 0 13 10 0 0 4
738 196
741 196
741 138
184 138
7 2 14 0 0 12416 0 8 13 0 0 6
478 288
521 288
521 168
751 168
751 206
738 206
4 1 15 0 0 12416 0 13 8 0 0 6
738 226
742 226
742 277
541 277
541 228
478 228
3 5 16 0 0 20608 0 13 9 0 0 8
738 216
751 216
751 298
600 298
600 382
275 382
275 398
187 398
4 11 17 0 0 12416 0 9 11 0 0 4
187 388
245 388
245 423
725 423
3 10 18 0 0 12416 0 9 11 0 0 4
187 378
263 378
263 413
725 413
2 9 19 0 0 12416 0 9 11 0 0 4
187 368
289 368
289 403
725 403
7 1 2 0 0 0 0 9 7 0 0 3
187 418
231 418
231 466
8 1 20 0 0 4224 0 11 9 0 0 4
725 393
313 393
313 358
187 358
12 0 2 0 0 4096 0 11 0 0 29 2
725 433
670 433
7 0 2 0 0 0 0 11 0 0 29 2
725 383
670 383
6 0 2 0 0 0 0 11 0 0 29 2
725 373
670 373
1 1 2 0 0 8320 0 11 3 0 0 3
725 323
670 323
670 467
4 5 21 0 0 12416 0 10 11 0 0 4
184 128
332 128
332 363
725 363
4 3 22 0 0 4224 0 11 10 0 0 4
725 353
341 353
341 118
184 118
2 3 23 0 0 12416 0 10 11 0 0 4
184 108
350 108
350 343
725 343
1 2 24 0 0 12416 0 10 11 0 0 4
184 98
361 98
361 333
725 333
8 1 2 0 0 0 0 8 5 0 0 3
478 298
492 298
492 300
7 1 2 0 0 0 0 10 6 0 0 3
184 158
221 158
221 205
53
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 6
749 186 785 201
753 190 784 201
6 X REF+
-16 0 0 0 400 0 0 0 0 3 2 1 18
15 Times New Roman
0 0 0 43
771 474 972 524
775 478 970 516
43 TO MOTION INT.BOARD J4
PIN 7,8,32,33 resp.
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
41 563 153 587
45 567 149 583
13 TO Y AXIS 1CN
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 7
104 594 145 609
108 598 144 609
7 20 *PCO
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 6
103 583 141 598
107 587 140 598
6 19 PCO
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
44 480 156 504
48 484 152 500
13 TO X AXIS 1CN
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 7
105 510 146 525
109 514 145 525
7 25 *PCO
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 6
105 499 143 514
109 503 142 514
6 24 PCO
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
155 52 331 76
159 56 327 72
21 X AXIS 1CN(SGDA-04AS)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
120 316 304 340
124 320 300 336
22 Y AXIS 1CN(SGDB-15ADG)
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 10
95 170 143 185
99 174 142 185
10 13 +24V IN
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
133 53 157 77
137 57 153 73
2 TO
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
100 316 124 340
104 320 120 336
2 TO
-13 0 0 0 400 0 0 0 0 3 2 1 18
15 Times New Roman
0 0 0 30
796 179 882 236
800 183 881 228
30 TO I/O
INTERFACE 
BOARD  J11
-13 0 0 0 400 0 0 0 0 3 2 1 18
15 Times New Roman
0 0 0 44
793 345 888 420
797 349 887 409
44 TO MOTION
CONTROLLER
INTERFACE
BOARD  J13
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 10
101 430 149 445
105 433 148 444
10 47 +24V IN
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 7
101 420 141 435
105 424 140 435
7 40 S-ON
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 4
102 410 127 425
106 414 126 425
4 1 SG
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 5
102 400 132 415
106 404 131 415
5 10 SG
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 7
102 390 142 405
106 394 141 405
7 9 T-REF
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 7
103 381 144 396
107 385 143 396
7 34 *PAO
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 6
103 369 141 384
107 373 140 384
6 33 PAO
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 7
102 359 143 374
106 363 142 374
7 36 *PBO
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 6
103 349 141 364
107 353 140 364
6 35 PBO
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 7
95 159 135 174
99 163 134 174
7 14 S-ON
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 5
95 150 125 165
99 154 124 165
5 19 SG
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 4
96 140 121 155
100 144 120 155
4 2 SG
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 7
96 130 136 145
100 134 135 145
7 1 T-REF
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 7
96 120 137 135
100 124 136 135
7 21 *PAO
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 6
95 110 133 125
99 114 132 125
6 20 PAO
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 7
96 100 137 115
100 104 136 115
7 23 *PBO
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 6
96 89 134 104
100 93 133 104
6 22 PBO
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 3
755 415 776 430
759 419 775 430
3 *YB
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 2
754 406 772 421
758 410 771 421
2 YB
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 3
754 395 775 410
758 399 774 410
3 *YA
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 2
754 385 772 400
758 389 771 400
2 YA
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 3
754 425 780 440
758 429 779 440
3 GND
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 3
754 376 780 391
758 380 779 391
3 GND
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 3
754 366 780 381
758 370 779 381
3 GND
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 3
755 356 776 371
759 360 775 371
3 *XB
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 2
755 345 773 360
759 349 772 360
2 XB
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 3
754 335 775 350
758 339 774 350
3 *XA
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 2
755 326 773 341
759 329 772 340
2 XA
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 3
755 314 781 329
759 318 780 329
3 GND
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
587 223 643 247
591 227 639 243
6 Y REF-
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
579 189 635 213
583 193 631 209
6 X REF-
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
630 205 662 229
634 209 658 225
3 GND
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
644 179 676 203
648 183 672 199
3 GND
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 5
749 217 778 232
753 221 777 232
5 Y INH
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 6
748 207 784 222
752 211 783 222
6 Y REF+
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 5
749 196 778 211
753 200 777 211
5 X INH
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
717 97 749 121
721 101 745 117
3 GND
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
716 86 756 110
720 90 752 106
4 +24V
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
