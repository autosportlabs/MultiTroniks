CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
20 78 780 559
7 5.000 V
7 5.000 V
3 GND
1000 10
24 100 0 1 0
20 Package,Description,
61 C:\PROGRAM FILES\MICROCODE ENGINEERING\CIRCUITMAKER 6\BOM.DAT
0 7
20 78 780 559
143654930 0
0
0
0
0
0
0
40
10 TER BLOCK~
94 482 43 0 2 5
0 8 9
10 TER BLOCK~
1 0 0 0
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
8953 0 0
0
0
10 TER BLOCK~
94 482 53 0 2 5
0 8 10
10 TER BLOCK~
2 0 0 0
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
4441 0 0
0
0
10 TER BLOCK~
94 482 63 0 2 5
0 7 11
10 TER BLOCK~
3 0 0 0
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
3618 0 0
0
0
10 TER BLOCK~
94 482 73 0 2 5
0 7 12
10 TER BLOCK~
4 0 0 0
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
6153 0 0
0
0
10 TER BLOCK~
94 482 83 0 2 5
0 6 13
10 TER BLOCK~
5 0 0 0
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
5394 0 0
0
0
10 TER BLOCK~
94 482 93 0 2 5
0 6 14
10 TER BLOCK~
6 0 0 0
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
7734 0 0
0
0
10 TER BLOCK~
94 482 191 0 2 5
0 2 15
10 TER BLOCK~
7 0 0 0
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
9914 0 0
0
0
10 TER BLOCK~
94 482 201 0 2 5
0 16 17
10 TER BLOCK~
8 0 0 0
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
3747 0 0
0
0
10 TER BLOCK~
94 482 211 0 2 5
0 18 19
10 TER BLOCK~
9 0 0 0
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
3549 0 0
0
0
10 TER BLOCK~
94 482 221 0 2 5
0 20 21
10 TER BLOCK~
10 0 0 0
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
7931 0 0
0
0
10 TER BLOCK~
94 482 231 0 2 5
0 22 23
10 TER BLOCK~
11 0 0 0
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
9325 0 0
0
0
10 TER BLOCK~
94 482 241 0 2 5
0 24 25
10 TER BLOCK~
12 0 0 0
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
8903 0 0
0
0
10 TER BLOCK~
94 482 251 0 2 5
0 26 27
10 TER BLOCK~
13 0 0 0
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
3834 0 0
0
0
10 TER BLOCK~
94 482 261 0 2 5
0 28 29
10 TER BLOCK~
14 0 0 0
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
3363 0 0
0
0
10 TER BLOCK~
94 482 271 0 2 5
0 30 31
10 TER BLOCK~
15 0 0 0
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
7668 0 0
0
0
10 TER BLOCK~
94 482 281 0 2 5
0 3 32
10 TER BLOCK~
16 0 0 0
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
4718 0 0
0
0
10 TER BLOCK~
94 482 391 0 2 5
0 33 34
10 TER BLOCK~
17 0 0 0
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
3874 0 0
0
0
10 TER BLOCK~
94 482 401 0 2 5
0 35 36
10 TER BLOCK~
18 0 0 0
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
6671 0 0
0
0
10 TER BLOCK~
94 482 411 0 2 5
0 37 38
10 TER BLOCK~
19 0 0 0
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
3789 0 0
0
0
10 TER BLOCK~
94 482 421 0 2 5
0 39 40
10 TER BLOCK~
20 0 0 0
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
4871 0 0
0
0
10 TER BLOCK~
94 482 431 0 2 5
0 41 42
10 TER BLOCK~
21 0 0 0
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
3750 0 0
0
0
10 TER BLOCK~
94 482 441 0 2 5
0 5 43
10 TER BLOCK~
22 0 0 0
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
8778 0 0
0
0
10 TER BLOCK~
94 482 451 0 2 5
0 44 45
10 TER BLOCK~
23 0 0 0
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
538 0 0
0
0
10 TER BLOCK~
94 482 461 0 2 5
0 46 47
10 TER BLOCK~
24 0 0 0
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
6843 0 0
0
0
10 TER BLOCK~
94 482 471 0 2 5
0 48 49
10 TER BLOCK~
25 0 0 0
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
3136 0 0
0
0
10 TER BLOCK~
94 482 481 0 2 5
0 50 51
10 TER BLOCK~
26 0 0 0
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
5950 0 0
0
0
10 TER BLOCK~
94 482 291 0 2 5
0 52 53
10 TER BLOCK~
27 0 0 0
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
5670 0 0
0
0
10 TER BLOCK~
94 482 311 0 2 5
0 54 55
10 TER BLOCK~
28 0 0 0
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
6828 0 0
0
0
10 TER BLOCK~
94 482 301 0 2 5
0 56 57
10 TER BLOCK~
29 0 0 0
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
6735 0 0
0
0
10 TER BLOCK~
94 482 321 0 2 5
0 4 58
10 TER BLOCK~
30 0 0 0
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
8365 0 0
0
0
10 TER BLOCK~
94 482 331 0 2 5
0 59 60
10 TER BLOCK~
31 0 0 0
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
4132 0 0
0
0
10 TER BLOCK~
94 482 341 0 2 5
0 61 62
10 TER BLOCK~
32 0 0 0
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
4551 0 0
0
0
10 TER BLOCK~
94 482 351 0 2 5
0 63 64
10 TER BLOCK~
33 0 0 0
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
3635 0 0
0
0
10 TER BLOCK~
94 482 361 0 2 5
0 65 66
10 TER BLOCK~
34 0 0 0
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
3973 0 0
0
0
10 TER BLOCK~
94 482 371 0 2 5
0 67 68
10 TER BLOCK~
35 0 0 0
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
3851 0 0
0
0
10 TER BLOCK~
94 482 381 0 2 5
0 69 70
10 TER BLOCK~
36 0 0 0
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
8383 0 0
0
0
2 PS
94 153 71 0 5 11
0 71 72 8 5 2
2 PS
37 0 4480 512
6 24V/5A
-25 -4 17 4
2 PS
-7 -60 7 -52
0
0
0
0
0
0
11

0 2 3 1 4 5 2 3 1 4
5 0
0 0 0 512 1 0 0 0
2 PS
9334 0 0
0
0
2 PS
94 152 204 0 5 11
0 7 6 8 5 3
2 PS
38 0 4480 512
6 12V/5A
-27 -4 15 4
2 PS
-7 -60 7 -52
0
0
0
0
0
0
11

0 2 3 1 4 5 2 3 1 4
5 0
0 0 0 0 1 0 0 0
2 PS
7471 0 0
0
0
2 PS
94 152 349 0 5 11
0 7 6 8 5 4
2 PS
39 0 4480 512
6 5V/10A
-28 -5 14 3
2 PS
-7 -60 7 -52
0
0
0
0
0
0
11

0 2 3 1 4 5 2 3 1 4
5 0
0 0 0 0 1 0 0 0
2 PS
3334 0 0
0
0
2 PS
94 151 484 0 5 11
0 7 6 8 5 73
2 PS
40 0 4480 512
7 24V/16A
-30 -2 19 6
2 PS
-7 -60 7 -52
0
0
0
0
0
0
11

0 2 3 1 4 5 2 3 1 4
5 0
0 0 0 512 1 0 0 0
2 PS
3559 0 0
0
0
22
1 0 0 0 0 0 0 37 0 0 16 3
215 51
251 51
251 62
0 2 0 0 0 0 0 0 37 13 0 4
262 82
229 82
229 61
215 61
1 5 2 0 0 4224 0 7 37 0 0 4
464 190
283 190
283 101
214 101
5 1 3 0 0 12416 0 38 16 0 0 4
213 234
284 234
284 280
464 280
5 1 4 0 0 12416 0 39 30 0 0 4
213 379
283 379
283 320
464 320
4 0 5 0 0 4096 0 39 0 0 8 2
213 369
273 369
4 0 5 0 0 0 0 38 0 0 8 2
213 224
273 224
0 4 5 0 0 8320 0 0 37 9 0 3
273 440
273 91
214 91
4 1 5 0 0 0 0 40 22 0 0 4
212 504
273 504
273 440
464 440
2 0 6 0 0 4096 0 39 0 0 13 2
214 339
262 339
2 0 6 0 0 0 0 38 0 0 13 2
214 194
262 194
0 1 6 0 0 0 0 0 6 13 0 3
446 82
446 92
464 92
2 1 6 0 0 8320 0 40 5 0 0 4
213 474
262 474
262 82
464 82
0 1 7 0 0 4096 0 0 40 15 0 3
251 329
251 464
213 464
0 1 7 0 0 4096 0 0 39 16 0 3
251 184
251 329
214 329
0 1 7 0 0 4224 0 0 38 17 0 4
445 62
251 62
251 184
214 184
1 1 7 0 0 0 0 3 4 0 0 4
464 62
445 62
445 72
464 72
3 0 8 0 0 4096 0 38 0 0 20 2
214 174
239 174
3 0 8 0 0 0 0 39 0 0 20 2
214 319
239 319
0 3 8 0 0 4224 0 0 40 22 0 3
239 41
239 454
213 454
1 0 8 0 0 0 0 2 0 0 22 3
464 52
445 52
445 41
1 3 8 0 0 0 0 1 37 0 0 3
464 42
464 41
215 41
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
