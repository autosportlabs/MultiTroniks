CircuitMaker Text
5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 25 3
0 66 799 572
7 5.000 V
7 5.000 V
3 GND
0 66 799 572
145752082 0
0
0
0
0
0
0
38
7 Ground~
168 833 1202 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8953 0 0
0
0
7 Ground~
168 403 1228 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4441 0 0
0
0
7 Ground~
168 82 1137 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3618 0 0
0
0
7 Ground~
168 1909 676 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6153 0 0
0
0
7 Ground~
168 1630 629 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5394 0 0
0
0
7 Ground~
168 1354 331 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7734 0 0
0
0
7 Ground~
168 804 596 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9914 0 0
0
0
7 Ground~
168 544 575 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3747 0 0
0
0
7 Ground~
168 743 287 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3549 0 0
0
0
7 Ground~
168 217 215 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7931 0 0
0
0
7 Ground~
168 271 347 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9325 0 0
0
0
7 Ground~
168 159 695 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8903 0 0
0
0
7 Ground~
168 1310 685 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3834 0 0
0
0
5 SIP8~
219 1731 491 0 8 17
0 22 20 166 167 168 21 19 169
0
0 0 608 90
4 CONN
9 2 37 10
2 J7
-9 -20 5 -12
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 512 1 0 0 0
1 J
3363 0 0
0
0
5 SIP8~
219 742 256 0 8 17
0 42 40 170 171 2 41 39 172
0
0 0 608 90
4 CONN
9 2 37 10
2 J6
-12 -20 2 -12
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 512 1 0 0 0
1 J
7668 0 0
0
0
5 CON50
94 967 497 0 101 101
0 2 173 34 33 32 31 174 175 176
177 178 179 61 180 181 182 88 183 184
185 90 89 186 187 2 188 2 38 37
36 35 189 190 191 2 192 193 58 194
195 196 85 197 198 199 87 86 200 201
2 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 -1610612324
5 CON50
145 0 2560 0
5 CON50
-18 -132 17 -124
2 J2
-8 -142 6 -134
0
0
0
0
0
0
101

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 21 22 23 24 25 26 27 28 29
30 31 32 33 34 35 36 37 38 39
40 41 42 43 44 45 46 47 48 49
50 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 21 22 23 24 25 26 27 28 29
30 31 32 33 34 35 36 37 38 39
40 41 42 43 44 45 46 47 48 49
50 0
0 0 0 512 1 0 0 0
1 J
4718 0 0
0
0
5 DB-37
94 106 495 0 75 75
0 2 70 71 37 35 33 31 45 43
68 41 39 202 119 117 115 72 47 2
2 70 38 36 34 32 46 44 42 40
203 120 118 116 114 69 2 47 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 -1610612428
5 DB-37
146 0 2688 512
4 DB37
-14 -200 14 -192
2 P1
-8 -201 6 -193
0
0
0
0
0
5 DB37M
75

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 21 22 23 24 25 26 27 29 30
31 32 33 34 35 28 37 36 1 2
3 4 5 6 7 8 9 10 11 12
13 14 15 16 17 18 19 20 21 22
23 24 25 26 27 29 30 31 32 33
34 35 28 37 36 0
0 0 0 512 1 0 0 0
1 J
3874 0 0
0
0
5 DB-37
94 1255 482 0 75 75
0 2 70 241 242 29 27 62 25 23
65 21 19 243 112 110 244 107 47 2
2 70 245 30 28 63 26 24 22 20
246 113 111 247 109 66 2 47 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 -1610612428
5 DB-37
147 0 2688 512
4 DB37
-14 -200 14 -192
2 P2
-7 -210 7 -202
0
0
0
0
0
5 DB37M
75

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 21 22 23 24 25 26 27 29 30
31 32 33 34 35 28 37 36 1 2
3 4 5 6 7 8 9 10 11 12
13 14 15 16 17 18 19 20 21 22
23 24 25 26 27 29 30 31 32 33
34 35 28 37 36 0
0 0 0 512 1 0 0 0
1 J
6671 0 0
0
0
5 CON50
94 1634 471 0 101 101
0 285 2 26 25 24 23 286 287 288
289 290 291 64 292 293 294 76 295 296
297 78 77 298 299 2 300 2 22 21
20 19 301 302 303 2 304 305 306 307
308 309 73 310 311 312 75 74 313 314
2 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 -1610612324
5 CON50
148 0 2688 0
5 CON50
-18 -132 17 -124
2 J3
-8 -142 6 -134
0
0
0
0
0
0
101

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 21 22 23 24 25 26 27 28 29
30 31 32 33 34 35 36 37 38 39
40 41 42 43 44 45 46 47 48 49
50 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 21 22 23 24 25 26 27 28 29
30 31 32 33 34 35 36 37 38 39
40 41 42 43 44 45 46 47 48 49
50 0
0 0 0 512 1 0 0 0
1 J
3789 0 0
0
0
5 CON50
94 649 502 0 101 101
0 315 2 46 45 44 43 316 317 318
319 320 321 67 322 323 324 82 325 326
327 84 83 328 329 2 330 2 42 41
40 39 331 332 333 2 334 335 336 337
338 339 79 340 341 342 81 80 343 344
2 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 -1610612476
5 CON50
149 0 2560 0
5 CON50
-18 -132 17 -124
2 J1
-8 -142 6 -134
0
0
0
0
0
0
101

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 21 22 23 24 25 26 27 28 29
30 31 32 33 34 35 36 37 38 39
40 41 42 43 44 45 46 47 48 49
50 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 21 22 23 24 25 26 27 28 29
30 31 32 33 34 35 36 37 38 39
40 41 42 43 44 45 46 47 48 49
50 0
0 0 0 512 1 0 0 0
1 J
4871 0 0
0
0
5 DB-37
94 36 939 0 75 75
0 345 346 111 113 120 117 118 7 9
110 2 347 2 348 2 349 2 350 2
351 352 353 354 355 109 6 8 114 112
119 115 116 11 12 10 14 13 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 -1610612428
5 DB-37
150 0 2560 512
4 DB37
-14 -200 14 -192
5 P1DIO
-24 208 11 216
0
0
0
0
0
5 DB37M
75

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 21 22 23 24 25 26 27 29 30
31 32 33 34 35 28 37 36 1 2
3 4 5 6 7 8 9 10 11 12
13 14 15 16 17 18 19 20 21 22
23 24 25 26 27 29 30 31 32 33
34 35 28 37 36 0
0 0 0 512 1 0 0 0
1 J
3750 0 0
0
0
5 CON50
94 1947 488 0 101 101
0 393 2 100 99 98 97 51 50 394
395 396 397 61 398 399 400 93 401 402
403 92 91 404 405 2 406 2 18 17
16 15 49 48 407 2 408 409 58 410
411 412 96 413 414 415 95 94 416 417
2 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 -1610612324
5 CON50
151 0 2688 0
5 CON50
-18 -132 17 -124
2 J4
-8 -142 6 -134
0
0
0
0
0
0
101

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 21 22 23 24 25 26 27 28 29
30 31 32 33 34 35 36 37 38 39
40 41 42 43 44 45 46 47 48 49
50 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 21 22 23 24 25 26 27 28 29
30 31 32 33 34 35 36 37 38 39
40 41 42 43 44 45 46 47 48 49
50 0
0 0 0 512 1 0 0 0
1 J
8778 0 0
0
0
5 CON10
94 736 848 0 10 21
0 418 107 59 105 102 419 108 60 106
103
5 CON10
152 0 4608 0
0
2 J5
-17 -61 -3 -53
0
0
0
0
0
5 IDC10
21

0 2 4 6 8 10 1 3 5 7
9 2 4 6 8 10 1 3 5 7
9 0
0 0 0 512 1 0 0 0
1 A
538 0 0
0
0
5 CON10
94 752 1207 0 10 21
0 2 2 108 3 4 2 2 72 5
3
5 CON10
153 0 4608 0
0
5 J3DIO
-27 -60 8 -52
0
0
0
0
0
5 IDC10
21

0 2 4 6 8 10 1 3 5 7
9 2 4 6 8 10 1 3 5 7
9 0
0 0 0 0 1 0 0 0
1 A
6843 0 0
0
0
5 CON10
94 1952 861 0 10 21
0 92 93 95 96 420 421 91 422 94
423
5 CON10
154 0 4608 0
0
6 J11DIO
-32 -60 10 -52
0
0
0
0
0
5 IDC10
21

0 2 4 6 8 10 1 3 5 7
9 2 4 6 8 10 1 3 5 7
9 0
0 0 0 512 1 0 0 0
1 A
3136 0 0
0
0
5 CON10
94 989 278 0 10 21
0 90 88 87 85 424 425 89 426 86
427
5 CON10
155 0 4608 0
0
3 J10
-22 15 -1 23
0
0
0
0
0
5 IDC10
21

0 2 4 6 8 10 1 3 5 7
9 2 4 6 8 10 1 3 5 7
9 0
0 0 0 512 1 0 0 0
1 A
5950 0 0
0
0
5 CON20
94 1480 194 0 20 41
0 428 83 429 80 430 77 431 74 432
433 84 82 81 79 78 76 75 73 434
435
5 CON20
156 0 4608 0
0
3 J11
-8 -66 13 -58
0
0
0
0
0
0
41

0 1 3 5 7 9 11 13 15 17
19 2 4 6 8 10 12 14 16 18
20 1 3 5 7 9 11 13 15 17
19 2 4 6 8 10 12 14 16 18
20 0
0 0 0 512 1 0 0 0
1 J
5670 0 0
0
0
4 CON4
94 192 147 0 4 9
0 47 70 71 2
4 CON4
157 0 4608 0
4 CON4
-16 -36 12 -28
2 J8
-11 -42 3 -34
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
1 J
6828 0 0
0
0
4 TER3
94 1729 352 0 3 7
0 30 100 55
4 TER3
158 0 0 512
0
0
0
0
0
0
0
0
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 J
6735 0 0
0
0
4 TER3
94 1799 376 0 3 7
0 29 99 54
4 TER3
159 0 0 512
0
0
0
0
0
0
0
0
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 J
8365 0 0
0
0
4 TER3
94 1732 421 0 3 7
0 28 98 53
4 TER3
160 0 0 512
0
0
0
0
0
0
0
0
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 J
4132 0 0
0
0
4 TER3
94 1832 319 0 3 7
0 27 97 52
4 TER3
161 0 0 512
0
0
0
0
0
0
0
0
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 J
4551 0 0
0
0
4 TER3
94 827 794 0 3 7
0 57 18 106
4 TER3
162 0 0 270
0
0
0
0
0
0
0
0
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 J
3635 0 0
0
0
4 TER3
94 857 871 0 3 7
0 104 17 105
4 TER3
163 0 0 270
0
0
0
0
0
0
0
0
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 J
3973 0 0
0
0
4 TER3
94 901 899 0 3 7
0 56 16 103
4 TER3
164 0 0 270
0
0
0
0
0
0
0
0
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 J
3851 0 0
0
0
4 TER3
94 967 895 0 3 7
0 101 15 102
4 TER3
165 0 0 270
0
0
0
0
0
0
0
0
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 J
8383 0 0
0
0
5 CON20
94 1095 838 0 20 41
0 531 54 52 532 104 101 51 49 533
47 55 53 534 57 56 535 50 48 536
47
5 CON20
166 0 4608 0
0
3 J13
-11 -66 10 -58
0
0
0
0
0
0
41

0 1 3 5 7 9 11 13 15 17
19 2 4 6 8 10 12 14 16 18
20 1 3 5 7 9 11 13 15 17
19 2 4 6 8 10 12 14 16 18
20 0
0 0 0 512 1 0 0 0
1 J
9334 0 0
0
0
5 CON62
94 519 1331 0 125 125
0 2 70 69 68 67 46 45 44 43
42 41 40 39 38 37 36 35 34 33
32 31 552 6 7 8 9 10 11 12
13 14 553 554 555 4 3 5 15 16
17 18 19 20 21 22 23 24 25 26
27 28 29 30 58 59 60 61 62 63
64 65 66 556 557 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 -1610612228
5 CON62
167 0 2176 0
0
0
0
0
0
0
0
0
125

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 21 22 23 24 25 26 27 28 29
30 31 32 33 34 35 36 37 38 39
40 41 42 43 44 45 46 47 48 49
50 51 52 53 54 55 56 57 58 59
60 61 62 63 64 1 2 3 4 5
6 7 8 9 10 11 12 13 14 15
16 17 18 19 20 21 22 23 24 25
26 27 28 29 30 31 32 33 34 35
36 37 38 39 40 41 42 43 44 45
46 47 48 49 50 51 52 53 54 55
56 57 58 59 60 0
0 0 0 0 1 1 0 0
1 J
7471 0 0
0
0
210
4 0 3 0 0 0 0 24 0 0 7 4
775 1197
801 1197
801 1255
686 1255
1 0 2 0 0 0 0 1 0 0 5 2
833 1196
833 1177
6 0 2 0 0 0 0 24 0 0 5 2
710 1167
695 1167
1 0 2 0 0 0 0 24 0 0 5 2
775 1167
833 1167
7 2 2 0 0 0 0 24 24 0 0 6
710 1177
695 1177
695 1145
833 1145
833 1177
775 1177
5 35 4 0 0 0 0 24 38 0 0 4
775 1207
782 1207
782 1444
551 1444
36 10 3 0 0 0 0 38 24 0 0 4
551 1435
686 1435
686 1207
710 1207
9 37 5 0 0 0 0 24 38 0 0 4
710 1197
674 1197
674 1426
551 1426
23 26 6 0 0 0 0 38 21 0 0 4
487 1399
95 1399
95 991
59 991
8 24 7 0 0 0 0 21 38 0 0 4
59 981
105 981
105 1408
487 1408
25 27 8 0 0 0 0 38 21 0 0 4
487 1417
114 1417
114 971
59 971
9 26 9 0 0 0 0 21 38 0 0 4
59 961
122 961
122 1426
487 1426
27 35 10 0 0 0 0 38 21 0 0 4
487 1435
131 1435
131 951
59 951
28 33 11 0 0 0 0 38 21 0 0 4
487 1444
141 1444
141 831
59 831
34 29 12 0 0 0 0 21 38 0 0 4
59 811
150 811
150 1453
487 1453
30 37 13 0 0 0 0 38 21 0 0 4
487 1462
160 1462
160 791
59 791
36 31 14 0 0 0 0 21 38 0 0 4
59 771
171 771
171 1471
487 1471
1 1 2 0 0 0 0 2 38 0 0 3
403 1222
403 1201
487 1201
0 38 15 0 0 0 0 0 38 167 0 3
1234 760
1234 1417
551 1417
0 39 16 0 0 0 0 0 38 170 0 3
1226 748
1226 1408
551 1408
0 40 17 0 0 0 0 0 38 172 0 3
1215 738
1215 1399
551 1399
0 41 18 0 0 0 0 0 38 175 0 3
1205 727
1205 1390
551 1390
42 0 19 0 0 0 0 38 0 0 184 3
551 1381
1474 1381
1474 645
0 43 20 0 0 0 0 0 38 185 0 3
1485 654
1485 1372
551 1372
44 0 21 0 0 0 0 38 0 0 186 3
551 1363
1495 1363
1495 665
0 45 22 0 0 0 0 0 38 187 0 3
1505 673
1505 1354
551 1354
46 0 23 0 0 0 0 38 0 0 188 4
551 1345
1514 1345
1514 504
1512 504
0 47 24 0 0 0 0 0 38 189 0 3
1522 514
1522 1336
551 1336
48 0 25 0 0 0 0 38 0 0 190 3
551 1327
1561 1327
1561 524
0 49 26 0 0 0 0 0 38 191 0 3
1551 534
1551 1318
551 1318
50 0 27 0 0 0 0 38 0 0 148 3
551 1309
1406 1309
1406 564
0 51 28 0 0 0 0 0 38 150 0 3
1396 574
1396 1300
551 1300
52 0 29 0 0 0 0 38 0 0 152 3
551 1291
1386 1291
1386 584
0 53 30 0 0 0 0 0 38 154 0 3
1376 594
1376 1282
551 1282
21 0 31 0 0 0 0 38 0 0 155 3
487 1381
180 1381
180 557
0 20 32 0 0 0 0 0 38 156 0 3
190 567
190 1372
487 1372
19 0 33 0 0 0 0 38 0 0 157 3
487 1363
198 1363
198 577
0 18 34 0 0 0 0 0 38 158 0 3
208 587
208 1354
487 1354
17 0 35 0 0 0 0 38 0 0 207 3
487 1345
218 1345
218 597
0 16 36 0 0 0 0 0 38 208 0 3
228 607
228 1336
487 1336
15 0 37 0 0 0 0 38 0 0 209 3
487 1327
237 1327
237 617
0 14 38 0 0 0 0 0 38 210 0 3
246 627
246 1318
487 1318
13 0 39 0 0 0 0 38 0 0 199 3
487 1309
256 1309
256 457
0 12 40 0 0 0 0 0 38 200 0 3
265 467
265 1300
487 1300
11 0 41 0 0 0 0 38 0 0 201 3
487 1291
274 1291
274 476
0 10 42 0 0 0 0 0 38 202 0 3
283 486
283 1282
487 1282
9 0 43 0 0 0 0 38 0 0 203 3
487 1273
292 1273
292 516
0 8 44 0 0 0 0 0 38 204 0 3
301 526
301 1264
487 1264
7 0 45 0 0 0 0 38 0 0 205 3
487 1255
311 1255
311 536
0 6 46 0 0 0 0 0 38 206 0 3
321 547
321 1246
487 1246
0 0 47 0 0 0 0 0 0 52 93 3
1124 883
1174 883
1174 208
10 20 47 0 0 0 0 37 37 0 0 6
1073 882
1069 882
1069 897
1124 897
1124 882
1117 882
33 18 48 0 0 0 0 22 37 0 0 6
1979 538
2102 538
2102 916
1603 916
1603 862
1117 862
8 32 49 0 0 0 0 37 22 0 0 6
1073 862
1062 862
1062 906
2091 906
2091 547
1979 547
17 8 50 0 0 0 0 37 22 0 0 6
1117 852
1160 852
1160 928
1842 928
1842 448
1915 448
7 7 51 0 0 0 0 37 22 0 0 6
1073 852
1028 852
1028 991
1831 991
1831 439
1915 439
3 3 52 0 0 0 0 32 37 0 0 6
1838 329
1856 329
1856 977
1039 977
1039 812
1073 812
3 12 53 0 0 0 0 31 37 0 0 6
1738 431
1784 431
1784 965
1147 965
1147 802
1117 802
3 2 54 0 0 0 0 30 37 0 0 6
1805 386
1818 386
1818 953
1052 953
1052 802
1073 802
11 3 55 0 0 0 0 37 29 0 0 6
1117 792
1148 792
1148 717
1773 717
1773 362
1735 362
1 15 56 0 0 0 0 35 37 0 0 6
911 893
928 893
928 932
1134 932
1134 832
1117 832
1 14 57 0 0 0 0 33 37 0 0 5
837 788
837 769
1135 769
1135 822
1117 822
54 0 58 0 0 0 0 38 0 0 146 3
551 1273
1192 1273
1192 770
55 3 59 0 0 0 0 38 23 0 0 6
551 1264
663 1264
663 953
776 953
776 828
759 828
8 56 60 0 0 0 0 23 38 0 0 4
694 829
649 829
649 1255
551 1255
57 0 61 0 0 0 0 38 0 0 145 8
551 1246
1672 1246
1672 792
1800 792
1800 494
1975 494
1975 493
1875 493
7 58 62 0 0 0 0 18 38 0 0 4
1278 544
1353 544
1353 1237
551 1237
59 25 63 0 0 0 0 38 18 0 0 4
551 1228
1363 1228
1363 554
1278 554
13 60 64 0 0 0 0 19 38 0 0 6
1602 476
1588 476
1588 1119
605 1119
605 1219
551 1219
61 10 65 0 0 0 0 38 18 0 0 6
551 1210
593 1210
593 1109
1342 1109
1342 484
1278 484
35 62 66 0 0 0 0 18 38 0 0 6
1278 494
1324 494
1324 1097
583 1097
583 1201
551 1201
5 13 67 0 0 0 0 38 20 0 0 6
487 1237
450 1237
450 766
561 766
561 507
617 507
10 4 68 0 0 0 0 17 38 0 0 4
129 497
441 497
441 1228
487 1228
3 35 69 0 0 0 0 38 17 0 0 4
487 1219
431 1219
431 507
129 507
0 2 70 0 0 0 0 0 38 111 0 4
342 657
343 657
343 1210
487 1210
1 0 2 0 0 0 0 3 0 0 80 2
82 1131
82 921
17 0 2 0 0 0 0 21 0 0 80 2
59 801
82 801
15 0 2 0 0 0 0 21 0 0 80 2
59 841
82 841
13 0 2 0 0 0 0 21 0 0 80 2
59 881
82 881
11 19 2 0 0 0 0 21 21 0 0 4
59 921
82 921
82 761
59 761
1 0 2 0 0 0 0 4 0 0 84 2
1909 670
1909 632
0 50 2 0 0 0 0 0 22 83 0 4
1998 520
1996 520
1996 385
1979 385
0 35 2 0 0 0 0 0 22 84 0 3
1998 593
1998 520
1979 520
0 27 2 0 0 0 0 0 22 85 0 5
1898 600
1898 632
1998 632
1998 592
1979 592
2 25 2 0 0 0 0 22 22 0 0 4
1915 394
1898 394
1898 601
1915 601
1 0 2 0 0 0 0 5 0 0 89 2
1630 623
1630 610
0 50 2 0 0 0 0 0 19 88 0 3
1682 503
1682 368
1666 368
0 35 2 0 0 0 0 0 19 89 0 3
1682 575
1682 503
1666 503
0 27 2 0 0 0 0 0 19 90 0 5
1580 582
1580 610
1682 610
1682 575
1666 575
2 25 2 0 0 0 0 19 19 0 0 4
1602 377
1580 377
1580 584
1602 584
0 0 70 0 0 0 0 0 0 92 111 5
1304 635
1303 635
1303 219
342 219
342 141
2 21 70 0 0 0 0 18 18 0 0 4
1278 644
1304 644
1304 634
1278 634
0 0 47 0 0 0 0 0 0 94 113 4
1322 324
1323 324
1323 208
241 208
37 18 47 0 0 0 0 18 18 0 0 4
1278 334
1322 334
1322 324
1278 324
19 0 2 0 0 0 0 18 0 0 96 3
1278 304
1302 304
1302 314
36 1 2 0 0 0 0 18 6 0 0 3
1278 314
1354 314
1354 325
1 0 2 0 0 0 0 7 0 0 98 3
804 590
804 572
846 572
1 0 2 0 0 0 0 16 0 0 101 3
935 394
846 394
846 610
50 0 2 0 0 0 0 16 0 0 100 3
999 394
1015 394
1015 530
0 35 2 0 0 0 0 0 16 101 0 3
1015 602
1015 529
999 529
25 27 2 0 0 0 0 16 16 0 0 6
935 610
846 610
846 639
1015 639
1015 601
999 601
1 0 2 0 0 0 0 8 0 0 103 3
544 569
544 555
572 555
2 0 2 0 0 0 0 20 0 0 106 4
617 408
572 408
572 615
573 615
50 0 2 0 0 0 0 20 0 0 105 3
681 399
696 399
696 535
0 35 2 0 0 0 0 0 20 106 0 3
696 607
696 534
681 534
25 27 2 0 0 0 0 20 20 0 0 6
617 615
573 615
573 639
696 639
696 606
681 606
1 5 2 0 0 0 0 9 15 0 0 3
743 281
744 281
744 265
1 4 2 0 0 0 0 10 28 0 0 3
217 209
217 161
206 161
3 3 71 0 0 0 0 17 28 0 0 4
129 637
331 637
331 151
206 151
0 21 70 0 0 0 0 0 17 111 0 3
159 657
159 647
129 647
2 2 70 0 0 0 0 28 17 0 0 4
206 141
342 141
342 657
129 657
37 0 47 0 0 0 0 17 0 0 113 3
129 347
241 347
241 336
18 1 47 0 0 0 0 17 28 0 0 4
129 337
241 337
241 131
206 131
17 8 72 0 0 0 0 17 24 0 0 6
129 357
352 357
352 750
634 750
634 1188
710 1188
19 0 2 0 0 0 0 17 0 0 116 3
129 317
159 317
159 327
1 36 2 0 0 0 0 11 17 0 0 3
271 341
271 327
129 327
1 0 2 0 0 0 0 12 0 0 118 2
159 689
159 677
20 1 2 0 0 0 0 17 17 0 0 4
129 667
159 667
159 677
129 677
1 0 2 0 0 0 0 13 0 0 120 2
1310 679
1310 663
20 1 2 0 0 0 0 18 18 0 0 4
1278 654
1310 654
1310 664
1278 664
18 42 73 0 0 0 0 27 19 0 0 4
1502 218
1709 218
1709 440
1666 440
8 47 74 0 0 0 0 27 19 0 0 6
1458 218
1437 218
1437 270
1699 270
1699 395
1666 395
17 46 75 0 0 0 0 27 19 0 0 4
1502 208
1690 208
1690 404
1666 404
16 17 76 0 0 0 0 27 19 0 0 4
1502 198
1571 198
1571 512
1602 512
22 6 77 0 0 0 0 19 27 0 0 6
1602 557
1532 557
1532 258
1445 258
1445 198
1458 198
15 21 78 0 0 0 0 27 19 0 0 4
1502 188
1541 188
1541 548
1602 548
14 42 79 0 0 0 0 27 20 0 0 6
1502 178
1538 178
1538 88
807 88
807 471
681 471
4 47 80 0 0 0 0 27 20 0 0 4
1458 178
798 178
798 426
681 426
13 46 81 0 0 0 0 27 20 0 0 6
1502 168
1527 168
1527 98
789 98
789 435
681 435
17 12 82 0 0 0 0 20 27 0 0 6
617 543
580 543
580 110
1517 110
1517 158
1502 158
2 22 83 0 0 0 0 27 20 0 0 4
1458 158
589 158
589 588
617 588
21 11 84 0 0 0 0 20 27 0 0 6
617 579
599 579
599 119
1508 119
1508 148
1502 148
4 42 85 0 0 0 0 26 16 0 0 4
1012 268
1053 268
1053 466
999 466
9 47 86 0 0 0 0 26 16 0 0 6
947 268
910 268
910 325
1035 325
1035 421
999 421
3 46 87 0 0 0 0 26 16 0 0 4
1012 258
1044 258
1044 430
999 430
2 17 88 0 0 0 0 26 16 0 0 6
1012 248
1024 248
1024 297
856 297
856 538
935 538
7 22 89 0 0 0 0 26 16 0 0 4
947 248
865 248
865 583
935 583
1 21 90 0 0 0 0 26 16 0 0 6
1012 238
1034 238
1034 307
874 307
874 574
935 574
22 7 91 0 0 0 0 22 25 0 0 4
1915 574
1868 574
1868 831
1910 831
21 1 92 0 0 0 0 22 25 0 0 6
1915 565
1878 565
1878 800
1977 800
1977 821
1975 821
17 2 93 0 0 0 0 22 25 0 0 6
1915 529
1888 529
1888 792
1988 792
1988 831
1975 831
47 9 94 0 0 0 0 22 25 0 0 6
1979 412
2082 412
2082 782
1898 782
1898 851
1910 851
46 3 95 0 0 0 0 22 25 0 0 4
1979 421
2072 421
2072 841
1975 841
42 4 96 0 0 0 0 22 25 0 0 4
1979 457
2062 457
2062 851
1975 851
13 13 61 0 0 0 0 16 22 0 0 8
935 502
919 502
919 316
1112 316
1112 281
1875 281
1875 493
1915 493
38 38 58 0 0 0 0 22 16 0 0 6
1979 493
2049 493
2049 770
1192 770
1192 502
999 502
2 6 97 0 0 0 0 32 22 0 0 4
1838 319
1866 319
1866 430
1915 430
6 1 27 0 0 0 0 18 32 0 0 6
1278 564
1406 564
1406 290
1845 290
1845 309
1838 309
5 2 98 0 0 0 0 22 31 0 0 2
1915 421
1738 421
24 1 28 0 0 0 0 18 31 0 0 6
1278 574
1397 574
1397 300
1781 300
1781 411
1738 411
4 2 99 0 0 0 0 22 30 0 0 4
1915 412
1829 412
1829 376
1805 376
5 1 29 0 0 0 0 18 30 0 0 6
1278 584
1386 584
1386 311
1815 311
1815 366
1805 366
3 2 100 0 0 0 0 22 29 0 0 4
1915 403
1838 403
1838 352
1735 352
23 1 30 0 0 0 0 18 29 0 0 6
1278 594
1376 594
1376 322
1745 322
1745 342
1735 342
7 6 31 0 0 0 0 17 16 0 0 6
129 557
490 557
490 306
817 306
817 439
935 439
25 5 32 0 0 0 0 17 16 0 0 6
129 567
498 567
498 316
894 316
894 430
935 430
6 4 33 0 0 0 0 17 16 0 0 6
129 577
507 577
507 326
903 326
903 421
935 421
24 3 34 0 0 0 0 17 16 0 0 6
129 587
516 587
516 335
912 335
912 412
935 412
7 0 19 0 0 0 0 14 0 0 184 3
1751 500
1754 500
1754 539
6 0 21 0 0 0 0 14 0 0 186 4
1742 500
1743 500
1743 557
1744 557
2 0 20 0 0 0 0 14 0 0 185 4
1706 500
1706 533
1708 533
1708 548
1 0 22 0 0 0 0 14 0 0 187 4
1697 500
1698 500
1698 566
1699 566
0 7 39 0 0 0 0 0 15 199 0 3
739 570
762 570
762 265
0 6 41 0 0 0 0 0 15 201 0 3
719 589
753 589
753 265
0 2 40 0 0 0 0 0 15 200 0 4
715 579
715 564
717 564
717 265
0 1 42 0 0 0 0 0 15 202 0 4
706 597
706 582
708 582
708 265
2 31 15 0 0 0 0 36 22 0 0 5
967 889
967 760
2042 760
2042 556
1979 556
6 1 101 0 0 0 0 37 36 0 0 3
1073 842
977 842
977 889
3 5 102 0 0 0 0 36 23 0 0 3
957 889
957 848
759 848
2 30 16 0 0 0 0 35 22 0 0 5
901 893
901 748
2031 748
2031 565
1979 565
10 3 103 0 0 0 0 23 35 0 0 5
694 848
685 848
685 894
891 894
891 893
2 29 17 0 0 0 0 34 22 0 0 5
857 865
857 738
2022 738
2022 574
1979 574
1 5 104 0 0 0 0 34 37 0 0 3
867 865
867 832
1073 832
4 3 105 0 0 0 0 23 34 0 0 3
759 838
847 838
847 865
2 28 18 0 0 0 0 33 22 0 0 5
827 788
827 727
2010 727
2010 583
1979 583
9 3 106 0 0 0 0 23 33 0 0 5
694 838
659 838
659 751
817 751
817 788
2 17 107 0 0 0 0 23 18 0 0 6
759 818
798 818
798 707
1415 707
1415 344
1278 344
7 3 108 0 0 0 0 23 24 0 0 6
694 818
672 818
672 921
818 921
818 1187
775 1187
34 25 109 0 0 0 0 18 21 0 0 4
1278 354
1425 354
1425 1011
59 1011
15 10 110 0 0 0 0 18 21 0 0 4
1278 384
1435 384
1435 941
59 941
32 3 111 0 0 0 0 18 21 0 0 4
1278 394
1445 394
1445 1081
59 1081
14 29 112 0 0 0 0 18 21 0 0 5
1278 404
1455 404
1455 912
59 912
59 911
31 4 113 0 0 0 0 18 21 0 0 4
1278 414
1464 414
1464 1061
59 1061
12 31 19 0 0 0 0 18 19 0 0 6
1278 444
1474 444
1474 645
1754 645
1754 539
1666 539
29 30 20 0 0 0 0 18 19 0 0 6
1278 454
1485 454
1485 655
1708 655
1708 548
1666 548
11 29 21 0 0 0 0 18 19 0 0 6
1278 464
1495 464
1495 665
1744 665
1744 557
1666 557
28 28 22 0 0 0 0 18 19 0 0 6
1278 474
1505 474
1505 673
1699 673
1699 566
1666 566
9 6 23 0 0 0 0 18 19 0 0 4
1278 504
1514 504
1514 413
1602 413
27 5 24 0 0 0 0 18 19 0 0 4
1278 514
1523 514
1523 404
1602 404
8 4 25 0 0 0 0 18 19 0 0 4
1278 524
1561 524
1561 395
1602 395
26 3 26 0 0 0 0 18 19 0 0 4
1278 534
1551 534
1551 386
1602 386
34 28 114 0 0 0 0 17 21 0 0 4
129 367
421 367
421 931
59 931
16 31 115 0 0 0 0 17 21 0 0 4
129 377
411 377
411 871
59 871
33 32 116 0 0 0 0 17 21 0 0 4
129 387
402 387
402 851
59 851
6 15 117 0 0 0 0 21 17 0 0 4
59 1021
392 1021
392 397
129 397
32 7 118 0 0 0 0 17 21 0 0 4
129 407
382 407
382 1001
59 1001
30 14 119 0 0 0 0 21 17 0 0 4
59 891
372 891
372 417
129 417
31 5 120 0 0 0 0 17 21 0 0 4
129 427
362 427
362 1041
59 1041
12 31 39 0 0 0 0 17 20 0 0 6
129 457
451 457
451 707
739 707
739 570
681 570
29 30 40 0 0 0 0 17 20 0 0 6
129 467
461 467
461 697
728 697
728 579
681 579
11 29 41 0 0 0 0 17 20 0 0 8
129 477
274 477
274 476
471 476
471 689
719 689
719 588
681 588
28 28 42 0 0 0 0 17 20 0 0 8
129 487
283 487
283 486
480 486
480 680
706 680
706 597
681 597
9 6 43 0 0 0 0 17 20 0 0 6
129 517
292 517
292 516
551 516
551 444
617 444
27 5 44 0 0 0 0 17 20 0 0 6
129 527
301 527
301 526
542 526
542 435
617 435
8 4 45 0 0 0 0 17 20 0 0 6
129 537
311 537
311 536
533 536
533 426
617 426
26 3 46 0 0 0 0 17 20 0 0 4
129 547
524 547
524 417
617 417
5 31 35 0 0 0 0 17 16 0 0 6
129 597
511 597
511 671
1074 671
1074 565
999 565
23 30 36 0 0 0 0 17 16 0 0 6
129 607
521 607
521 660
1065 660
1065 574
999 574
4 29 37 0 0 0 0 17 16 0 0 6
129 617
531 617
531 649
1056 649
1056 583
999 583
22 28 38 0 0 0 0 17 16 0 0 6
129 627
503 627
503 717
1048 717
1048 592
999 592
12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
679 763 775 787
683 767 771 783
11 Y INTERFACE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
695 1127 807 1151
699 1131 803 1147
13 RELAY CONTROL
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
1902 322 1982 346
1906 326 1978 342
9 XY ROTARY
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1570 325 1610 349
1574 329 1606 345
4 Z2T2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
942 340 998 364
946 344 994 360
6 XY LIN
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
624 335 664 359
628 339 660 355
4 Z1T1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
1684 449 1772 473
1688 453 1768 469
10 LASER ENC2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
695 204 783 228
699 208 779 224
10 LASER ENC1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
967 769 1079 793
971 773 1075 789
13 AC MOTOR ENC.
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 19
1873 868 2033 892
1877 872 2029 888
19  MOTOR DRIVE RORARY
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 15
922 204 1050 228
926 208 1046 224
15 MOTOR DRIVE LIN
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
0 1153 104 1177
4 1157 100 1173
12 TO DIO BOARD
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
