CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
610 490 30 100 9
19 79 772 576
7 5.000 V
7 5.000 V
3 GND
1000 10
24 100 0 1 0
20 Package,Description,
65 C:\PROGRAM FILES\MICROCODE ENGINEERING\CIRCUITMAKER 6 PRO\BOM.DAT
0 7
19 79 772 576
143654930 0
0
0
0
0
0
0
74
2 +V
167 890 609 0 1 3
0 0
0
0 0 53600 0
3 +5V
-10 -14 11 -6
3 V10
-11 -32 10 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
8953 0 0
0
0
5 SIP4~
219 311 824 0 1 9
0 0
0
0 0 608 270
4 CONN
9 2 37 10
3 J16
20 0 41 8
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 -1610612604
0 0 0 0 1 0 0 0
1 J
4441 0 0
0
0
5 SIP4~
219 414 825 0 1 9
0 0
0
0 0 608 270
4 CONN
9 2 37 10
3 J17
20 0 41 8
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 -1610612604
0 0 0 0 1 0 0 0
1 J
3618 0 0
0
0
5 SIP3~
219 532 827 0 1 7
0 0
0
0 0 608 270
4 CONN
-13 -25 15 -17
3 J18
18 -1 39 7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 -1610612604
0 0 0 0 1 0 0 0
1 J
6153 0 0
0
0
5 SIP4~
219 632 826 0 1 9
0 0
0
0 0 608 270
4 CONN
9 2 37 10
3 J19
20 0 41 8
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 -1610612604
0 0 0 0 1 0 0 0
1 J
5394 0 0
0
0
5 SIP3~
219 733 828 0 1 7
0 0
0
0 0 608 270
4 CONN
-13 -25 15 -17
3 J20
18 -1 39 7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 -1610612604
0 0 0 0 1 0 0 0
1 J
7734 0 0
0
0
5 SIP4~
219 917 828 0 1 9
0 0
0
0 0 608 270
4 CONN
9 2 37 10
3 J21
20 0 41 8
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 -1610612604
0 0 0 0 1 0 0 0
1 J
9914 0 0
0
0
5 SIP3~
219 1007 829 0 1 7
0 0
0
0 0 608 270
4 CONN
-13 -25 15 -17
3 J22
18 -1 39 7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 -1610612604
0 0 0 0 1 0 0 0
1 J
3747 0 0
0
0
5 SIP4~
219 1094 827 0 1 9
0 0
0
0 0 608 270
4 CONN
9 2 37 10
3 J23
20 0 41 8
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 -1610612604
0 0 0 0 1 0 0 0
1 J
3549 0 0
0
0
5 SIP3~
219 1188 827 0 1 7
0 0
0
0 0 608 270
4 CONN
-13 -25 15 -17
3 J24
18 -1 39 7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 -1610612604
0 0 0 0 1 0 0 0
1 J
7931 0 0
0
0
5 SIP2~
219 1184 184 0 1 5
0 0
0
0 0 608 90
4 CONN
9 2 37 10
3 J14
-14 -19 7 -11
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 -1610612604
0 0 0 0 1 0 0 0
1 J
9325 0 0
0
0
5 SIP2~
219 1127 183 0 1 5
0 0
0
0 0 608 90
4 CONN
9 2 37 10
3 J13
-14 -19 7 -11
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 -1610612604
0 0 0 0 1 0 0 0
1 J
8903 0 0
0
0
5 SIP2~
219 1073 183 0 1 5
0 0
0
0 0 608 90
4 CONN
9 2 37 10
3 J12
-14 -19 7 -11
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 -1610612604
0 0 0 0 1 0 0 0
1 J
3834 0 0
0
0
5 SIP2~
219 1017 183 0 1 5
0 0
0
0 0 608 90
4 CONN
9 2 37 10
3 J11
-14 -19 7 -11
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 -1610612604
0 0 0 0 1 0 0 0
1 J
3363 0 0
0
0
5 SIP3~
219 931 183 0 1 7
0 0
0
0 0 608 90
4 CONN
-13 -25 15 -17
3 J15
-11 -20 10 -12
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 -1610612604
0 0 0 0 1 0 0 0
1 J
7668 0 0
0
0
5 SIP2~
219 757 167 0 1 5
0 0
0
0 0 608 90
4 CONN
9 2 37 10
3 J26
10 -7 31 1
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 -1610612604
0 0 0 0 1 0 0 0
1 J
4718 0 0
0
0
5 SIP2~
219 711 167 0 1 5
0 0
0
0 0 608 90
4 CONN
9 2 37 10
3 J25
-37 -7 -16 1
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 -1610612604
0 0 0 0 1 0 0 0
1 J
3874 0 0
0
0
5 SIP2~
219 620 167 0 1 5
0 0
0
0 0 608 90
4 CONN
9 2 37 10
3 J10
10 -7 31 1
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 -1610612604
0 0 0 0 1 0 0 0
1 J
6671 0 0
0
0
5 SIP2~
219 571 166 0 1 5
0 0
0
0 0 608 90
4 CONN
9 2 37 10
2 J9
-28 -6 -14 2
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 -1610612604
0 0 0 0 1 0 0 0
1 J
3789 0 0
0
0
5 SIP2~
219 496 165 0 1 5
0 0
0
0 0 608 90
4 CONN
9 2 37 10
2 J8
-29 -7 -15 1
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 -1610612604
0 0 0 0 1 0 0 0
1 J
4871 0 0
0
0
5 SIP2~
219 444 166 0 1 5
0 0
0
0 0 608 90
4 CONN
9 2 37 10
2 J7
-28 -6 -14 2
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 -1610612604
0 0 0 0 1 0 0 0
1 J
3750 0 0
0
0
5 SIP2~
219 389 166 0 1 5
0 0
0
0 0 608 90
4 CONN
9 2 37 10
2 J6
-28 -7 -14 1
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 -1610612604
0 0 0 0 1 0 0 0
1 J
8778 0 0
0
0
5 SIP2~
219 335 165 0 1 5
0 0
0
0 0 608 90
4 CONN
9 2 37 10
2 J5
-29 -6 -15 2
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 -1610612604
0 0 0 0 1 0 0 0
1 J
538 0 0
0
0
5 SIP2~
219 283 164 0 1 5
0 0
0
0 0 608 90
4 CONN
9 2 37 10
2 J4
-30 -7 -16 1
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 -1610612604
0 0 0 0 1 0 0 0
1 J
6843 0 0
0
0
5 SIP3~
219 177 164 0 1 7
0 0
0
0 0 608 90
4 CONN
-13 -25 15 -17
2 J3
-30 -9 -16 -1
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 -1610612604
0 0 0 0 1 0 0 0
1 J
3136 0 0
0
0
7 Ground~
168 1217 416 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5950 0 0
0
0
10 Capacitor~
219 1234 390 0 2 5
0 2 3
0
0 0 832 0
6 0.01uF
-21 -18 21 -10
2 C6
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 CAP0.2
5

0 1 2 1 2 -1610612703
67 0 0 0 1 0 0 0
1 C
5670 0 0
0
0
2 +V
167 1094 535 0 1 3
0 11
0
0 0 53728 0
2 5V
-7 -22 7 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6828 0 0
0
0
2 +V
167 1262 367 0 1 3
0 3
0
0 0 53600 0
3 +5V
-11 -14 10 -6
2 V2
-8 -24 6 -16
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6735 0 0
0
0
7 Ground~
168 1202 606 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8365 0 0
0
0
7 Ground~
168 1041 736 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4132 0 0
0
0
7 Ground~
168 998 401 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4551 0 0
0
0
7 Ground~
168 923 212 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3635 0 0
0
0
7 Ground~
168 869 252 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3973 0 0
0
0
7 Ground~
168 868 674 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3851 0 0
0
0
2 +V
167 124 182 0 1 3
0 36
0
0 0 53600 0
3 +5V
7 1 28 9
2 V3
10 -9 24 -1
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8383 0 0
0
0
7 Ground~
168 593 231 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9334 0 0
0
0
10 Capacitor~
219 593 213 0 2 5
0 2 37
0
0 0 832 90
6 0.01uF
-56 11 -14 19
2 C2
-42 1 -28 9
0
0
11 %D %1 %2 %V
0
0
6 CAP0.2
5

0 1 2 1 2 -1610612676
67 0 0 0 1 0 0 0
1 C
7471 0 0
0
0
7 Ground~
168 622 231 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3334 0 0
0
0
7 Ground~
168 619 527 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3559 0 0
0
0
10 Capacitor~
219 619 506 0 2 5
0 2 42
0
0 0 832 90
6 0.01uF
-43 -17 -1 -9
2 C4
-29 -27 -15 -19
0
0
11 %D %1 %2 %V
0
0
6 CAP0.2
5

0 1 2 1 2 -1610612720
67 0 0 0 1 0 0 0
1 C
984 0 0
0
0
2 +V
167 639 692 0 1 3
0 43
0
0 0 53600 0
3 +5V
-29 -4 -8 4
2 V4
-26 -14 -12 -6
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7557 0 0
0
0
2 +V
167 265 750 0 1 3
0 8
0
0 0 53600 0
3 +5V
-10 -14 11 -6
2 V5
-7 -24 7 -16
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3146 0 0
0
0
7 Ground~
168 224 831 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5687 0 0
0
0
7 Ground~
168 207 300 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7939 0 0
0
0
10 Polar Cap~
219 208 283 0 2 5
0 50 2
0
0 0 832 270
5 200uF
-16 -32 19 -24
2 C8
-6 -42 8 -34
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 -1610612720
67 0 0 0 1 0 0 0
1 C
3308 0 0
0
0
2 +V
167 250 264 0 1 3
0 50
0
0 0 53600 270
3 24V
0 -12 21 -4
2 V6
3 -22 17 -14
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3408 0 0
0
0
7 Ground~
168 205 666 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9773 0 0
0
0
10 Polar Cap~
219 206 639 0 2 5
0 51 2
0
0 0 832 270
5 200uF
10 5 45 13
2 C3
16 -4 30 4
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 -1610612676
67 0 0 0 1 0 0 0
1 C
691 0 0
0
0
7 Ground~
168 405 609 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7834 0 0
0
0
10 Capacitor~
219 405 590 0 2 5
0 2 52
0
0 0 832 90
6 0.01uF
-44 -12 -2 -4
2 C5
-23 -20 -9 -12
0
0
11 %D %1 %2 %V
0
0
6 CAP0.2
5

0 1 2 1 2 -1610612720
67 0 0 0 1 0 0 0
1 C
3588 0 0
0
0
7 Ground~
168 239 235 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4528 0 0
0
0
10 Capacitor~
219 239 219 0 2 5
0 2 50
0
0 0 832 90
5 0.1uF
-38 -13 -3 -5
2 C1
7 -14 21 -6
0
0
11 %D %1 %2 %V
0
0
6 CAP0.2
5

0 1 2 1 2 -1610612704
67 0 0 0 1 0 0 0
1 C
3303 0 0
0
0
7 Ground~
168 147 275 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9654 0 0
0
0
7 Ground~
168 329 389 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9791 0 0
0
0
2 +V
167 676 480 0 1 3
0 42
0
0 0 53600 0
3 +5V
-12 -13 9 -5
2 V7
-9 -23 5 -15
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4589 0 0
0
0
7 Ground~
168 640 667 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
964 0 0
0
0
7 Ground~
168 365 746 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9151 0 0
0
0
2 +V
167 449 557 0 1 3
0 52
0
0 0 53600 0
3 +5V
-14 -12 7 -4
2 V8
-11 -22 3 -14
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4745 0 0
0
0
2 +V
167 237 610 0 1 3
0 51
0
0 0 53600 270
3 +5V
2 -4 23 4
2 V9
5 -14 19 -6
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8433 0 0
0
0
7 Ground~
168 163 667 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4221 0 0
0
0
6 26LS31
94 411 684 0 16 33
0 81 79 72 87 74 73 80 2 48
76 75 2 78 77 49 52
6 26LS31
1 0 6400 0
6 26LS31
-20 -57 22 -49
0
0
0
0
0
0
5 DIP16
33

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 1 2 3
4 5 6 7 8 9 10 11 12 13
14 15 16 -1610612488
0 0 0 512 1 1 0 0
1 U
8348 0 0
0
0
5 CON34
94 140 475 0 34 69
0 2 2 51 51 37 39 79 72 73
74 75 76 77 78 71 70 69 68 67
66 65 64 63 62 61 60 59 58 35
41 50 50 2 2
5 CON34
2 0 4608 0
5 CON34
-20 -186 15 -178
2 J1
-8 -186 6 -178
0
0
0
0
0
5 SIP34
69

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 21 22 23 24 25 26 27 28 29
30 31 32 33 34 1 2 3 4 5
6 7 8 9 10 11 12 13 14 15
16 17 18 19 20 21 22 23 24 25
26 27 28 29 30 31 32 33 34 0
0 0 0 0 1 0 0 0
1 J
5299 0 0
0
0
6 26LS31
94 640 597 0 16 33
0 47 71 70 202 68 69 45 2 44
67 66 2 64 65 46 42
6 26LS31
4 0 6528 0
6 26LS31
-20 -56 22 -48
0
0
0
0
0
0
5 DIP16
33

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 1 2 3
4 5 6 7 8 9 10 11 12 13
14 15 16 -1610612720
0 0 0 512 1 1 0 0
1 U
7393 0 0
0
0
4 2003
94 373 335 0 16 33
0 237 58 59 60 61 62 63 2 238
38 57 56 55 54 53 50
4 2003
5 0 6784 0
2 IC
-8 -56 6 -48
2 U5
-6 -54 8 -46
0
0
0
0
0
0
33

0 1 2 3 4 5 6 7 8 16
15 14 13 12 11 10 9 1 2 3
4 5 6 7 8 16 15 14 13 12
11 10 9 0
0 0 0 512 1 1 0 0
1 U
6917 0 0
0
0
5 CON34
94 846 490 0 34 69
0 2 2 34 34 411 412 413 414 415
416 23 22 21 20 19 18 17 16 15
14 13 12 32 31 30 29 417 418 33
419 28 28 2 2
5 CON34
20 0 4608 0
5 CON34
-20 -186 15 -178
2 J2
-10 -186 4 -178
0
0
0
0
0
5 SIP34
69

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 21 22 23 24 25 26 27 28 29
30 31 32 33 34 1 2 3 4 5
6 7 8 9 10 11 12 13 14 15
16 17 18 19 20 21 22 23 24 25
26 27 28 29 30 31 32 33 34 0
0 0 0 512 1 0 0 0
1 J
8767 0 0
0
0
6 26LS31
94 1048 642 0 16 33
0 10 23 22 420 20 21 9 2 6
17 16 2 18 19 7 11
6 26LS31
21 0 6912 0
6 26LS31
-20 -56 22 -48
2 U3
-6 -66 8 -58
0
0
0
0
0
5 DIP16
33

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 1 2 3
4 5 6 7 8 9 10 11 12 13
14 15 16 -1610612487
0 0 0 512 1 1 0 0
1 U
3606 0 0
0
0
6 26LS31
94 1220 512 0 16 33
0 5 15 14 455 456 457 458 2 459
460 461 2 12 13 4 3
6 26LS31
22 0 6912 0
6 26LS31
-20 -56 22 -48
2 U4
-6 -66 8 -58
0
0
0
0
0
5 DIP16
33

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 1 2 3
4 5 6 7 8 9 10 11 12 13
14 15 16 -1610612488
0 0 0 512 1 1 0 0
1 U
6970 0 0
0
0
4 2003
94 1038 343 0 16 33
0 668 669 670 29 30 31 32 2 671
672 673 24 25 26 27 28
4 2003
32 0 6912 0
5 2003A
-18 -56 17 -48
2 U6
-8 -66 6 -58
0
0
0
0
0
0
33

0 1 2 3 4 5 6 7 8 16
15 14 13 12 11 10 9 1 2 3
4 5 6 7 8 16 15 14 13 12
11 10 9 0
0 0 0 512 1 1 0 0
1 U
343 0 0
0
0
9 Resistor~
219 124 220 0 4 5
0 35 36 0 1
0
0 0 864 90
2 1k
8 -5 22 3
2 R1
8 -15 22 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612712
82 0 0 0 1 0 0 0
1 R
7197 0 0
0
0
9 Resistor~
219 661 732 0 4 5
0 44 43 0 1
0
0 0 352 90
3 2K2
5 -5 26 3
3 R10
5 -15 26 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612676
82 0 0 0 1 0 0 0
1 R
3623 0 0
0
0
9 Resistor~
219 618 736 0 4 5
0 45 43 0 1
0
0 0 352 90
3 2K2
-26 -4 -5 4
3 R11
-26 -14 -5 -6
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612704
82 0 0 0 1 0 0 0
1 R
7656 0 0
0
0
9 Resistor~
219 312 608 0 4 5
0 81 52 0 1
0
0 0 864 90
3 2K2
1 17 22 25
2 R3
4 7 18 15
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612676
82 0 0 0 1 0 0 0
1 R
5365 0 0
0
0
9 Resistor~
219 338 610 0 4 5
0 80 52 0 1
0
0 0 864 90
3 2K2
3 -7 24 1
2 R4
6 -17 20 -9
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612704
82 0 0 0 1 0 0 0
1 R
4557 0 0
0
0
156
1 0 0 0 0 0 0 1 0 0 54 3
890 618
890 629
869 629
1 1 2 0 0 8192 0 27 26 0 0 3
1225 390
1217 390
1217 410
2 0 3 0 0 4096 0 27 0 0 18 2
1243 390
1262 390
15 2 4 0 0 16512 0 68 10 0 0 5
1252 486
1276 486
1276 629
1187 629
1187 819
1 1 5 0 0 8320 0 68 9 0 0 5
1188 476
1174 476
1174 771
1105 771
1105 819
9 2 6 0 0 8320 0 67 9 0 0 4
1080 676
1095 676
1095 819
1096 819
15 2 7 0 0 8320 0 67 8 0 0 5
1080 616
1119 616
1119 756
1006 756
1006 821
3 0 2 0 0 4096 0 7 0 0 11 2
910 820
910 799
1 0 2 0 0 4096 0 8 0 0 11 2
1015 821
1015 799
3 0 2 0 0 0 0 9 0 0 11 2
1087 819
1087 799
0 1 2 0 0 4096 0 0 10 87 0 3
741 799
1196 799
1196 819
4 0 8 0 0 4096 0 9 0 0 15 2
1078 819
1078 787
3 0 8 0 0 4096 0 8 0 0 15 2
997 821
997 787
4 0 8 0 0 0 0 7 0 0 15 2
901 820
901 787
0 3 8 0 0 4224 0 0 10 91 0 3
723 787
1178 787
1178 819
1 7 9 0 0 4224 0 7 67 0 0 3
928 820
928 666
1016 666
1 2 10 0 0 8320 0 67 7 0 0 3
1016 606
919 606
919 820
1 16 3 0 0 4224 0 29 68 0 0 3
1262 376
1262 476
1252 476
1 16 11 0 0 4224 0 28 67 0 0 3
1094 544
1094 606
1080 606
1 0 2 0 0 0 0 30 0 0 22 2
1202 600
1202 568
1 0 2 0 0 0 0 31 0 0 23 2
1041 730
1041 722
8 12 2 0 0 0 0 68 68 0 0 6
1188 546
1185 546
1185 568
1263 568
1263 516
1252 516
8 12 2 0 0 0 0 67 67 0 0 6
1016 676
1008 676
1008 722
1108 722
1108 646
1080 646
22 13 12 0 0 4224 0 66 68 0 0 4
860 444
1297 444
1297 506
1252 506
21 14 13 0 0 4224 0 66 68 0 0 4
860 454
1286 454
1286 496
1252 496
20 3 14 0 0 4224 0 66 68 0 0 4
860 464
1166 464
1166 496
1188 496
19 2 15 0 0 4224 0 66 68 0 0 4
860 474
1156 474
1156 486
1188 486
18 11 16 0 0 4224 0 66 67 0 0 4
860 484
1144 484
1144 656
1080 656
17 10 17 0 0 4224 0 66 67 0 0 4
860 494
1135 494
1135 666
1080 666
16 13 18 0 0 4224 0 66 67 0 0 4
860 504
1126 504
1126 636
1080 636
15 14 19 0 0 4224 0 66 67 0 0 4
860 514
1110 514
1110 626
1080 626
14 5 20 0 0 8320 0 66 67 0 0 4
860 524
931 524
931 646
1016 646
13 6 21 0 0 8320 0 66 67 0 0 4
860 534
944 534
944 656
1016 656
12 3 22 0 0 4224 0 66 67 0 0 4
860 544
957 544
957 626
1016 626
11 2 23 0 0 4224 0 66 67 0 0 4
860 553
967 553
967 616
1016 616
2 12 24 0 0 12416 0 14 69 0 0 5
1019 192
1019 241
1083 241
1083 337
1069 337
2 13 25 0 0 12416 0 13 69 0 0 5
1075 192
1075 226
1106 226
1106 347
1069 347
2 14 26 0 0 8320 0 12 69 0 0 4
1129 192
1128 192
1128 357
1069 357
2 15 27 0 0 4224 0 11 69 0 0 3
1186 193
1186 367
1069 367
16 0 28 0 0 8192 0 69 0 0 44 3
1069 377
1150 377
1150 213
1 0 28 0 0 0 0 14 0 0 44 2
1010 192
1010 213
1 0 28 0 0 0 0 13 0 0 44 2
1066 192
1066 213
1 0 28 0 0 0 0 12 0 0 44 2
1120 192
1120 213
0 1 28 0 0 4224 0 0 11 53 0 5
941 213
1150 213
1150 212
1177 212
1177 193
26 4 29 0 0 4224 0 66 69 0 0 4
860 404
953 404
953 337
1006 337
25 5 30 0 0 4224 0 66 69 0 0 4
860 414
963 414
963 347
1006 347
6 24 31 0 0 12416 0 69 66 0 0 4
1006 357
973 357
973 424
860 424
23 7 32 0 0 4224 0 66 69 0 0 4
860 434
986 434
986 367
1006 367
8 1 2 0 0 0 0 69 32 0 0 3
1006 377
998 377
998 395
29 2 33 0 0 8320 0 66 15 0 0 3
860 374
932 374
932 191
1 1 2 0 0 0 0 15 33 0 0 2
923 191
923 206
31 0 28 0 0 0 0 66 0 0 53 3
860 354
898 354
898 344
3 32 28 0 0 0 0 15 66 0 0 3
941 191
941 344
860 344
3 4 34 0 0 8320 0 66 66 0 0 4
860 634
869 634
869 624
860 624
1 0 2 0 0 0 0 66 0 0 56 2
860 654
868 654
2 1 2 0 0 0 0 66 35 0 0 3
860 644
868 644
868 668
34 0 2 0 0 0 0 66 0 0 58 2
860 324
898 324
1 33 2 0 0 0 0 34 66 0 0 5
869 246
869 237
898 237
898 334
860 334
1 0 35 0 0 8192 0 70 0 0 114 3
124 238
124 245
178 245
1 2 36 0 0 4224 0 36 70 0 0 2
124 191
124 202
1 1 2 0 0 0 0 38 37 0 0 2
593 222
593 225
2 0 37 0 0 4096 0 38 0 0 65 2
593 204
593 196
2 1 2 0 0 0 0 18 39 0 0 2
622 176
622 225
10 2 38 0 0 12416 0 65 19 0 0 5
404 309
465 309
465 212
573 212
573 175
0 1 37 0 0 4096 0 0 18 66 0 3
564 196
613 196
613 176
5 1 37 0 0 8320 0 63 19 0 0 7
154 599
247 599
247 298
317 298
317 269
564 269
564 175
2 6 39 0 0 8320 0 16 63 0 0 7
759 176
759 259
302 259
302 287
235 287
235 589
154 589
2 1 40 0 0 8320 0 17 16 0 0 4
713 176
713 201
750 201
750 176
30 1 41 0 0 20608 0 63 17 0 0 7
154 349
221 349
221 277
291 277
291 247
704 247
704 176
1 1 2 0 0 0 0 40 41 0 0 2
619 521
619 515
2 1 42 0 0 8192 0 41 56 0 0 3
619 497
619 489
676 489
1 0 43 0 0 4096 0 42 0 0 73 2
639 701
639 711
2 2 43 0 0 8320 0 72 71 0 0 4
618 718
618 711
661 711
661 714
1 0 44 0 0 4096 0 71 0 0 79 2
661 750
661 769
1 0 45 0 0 4096 0 72 0 0 78 2
618 754
618 769
0 1 8 0 0 0 0 0 43 91 0 3
295 787
265 787
265 759
15 2 46 0 0 8320 0 64 6 0 0 3
672 571
732 571
732 820
7 2 45 0 0 8320 0 64 5 0 0 5
608 621
586 621
586 769
634 769
634 818
9 1 44 0 0 8320 0 64 5 0 0 6
672 631
687 631
687 769
642 769
642 818
643 818
1 2 47 0 0 8320 0 64 4 0 0 3
608 561
531 561
531 819
9 2 48 0 0 16512 0 62 3 0 0 5
443 718
449 718
449 754
416 754
416 817
15 1 49 0 0 8320 0 62 3 0 0 5
443 658
484 658
484 765
425 765
425 817
3 0 2 0 0 0 0 5 0 0 87 2
625 818
625 799
1 0 2 0 0 0 0 4 0 0 87 2
540 819
540 799
3 0 2 0 0 0 0 3 0 0 87 2
407 817
407 799
3 0 2 0 0 0 0 2 0 0 87 2
304 816
304 799
1 1 2 0 0 8320 0 6 44 0 0 4
741 820
741 799
224 799
224 825
4 0 8 0 0 0 0 3 0 0 91 3
398 817
399 817
399 787
3 0 8 0 0 0 0 4 0 0 91 2
522 819
522 787
4 0 8 0 0 0 0 5 0 0 91 2
616 818
616 787
4 3 8 0 0 0 0 2 6 0 0 4
295 816
295 787
723 787
723 820
1 2 2 0 0 0 0 45 46 0 0 2
207 294
207 290
1 0 50 0 0 4096 0 46 0 0 95 2
207 273
207 263
16 0 50 0 0 8192 0 65 0 0 111 3
404 369
481 369
481 198
1 0 50 0 0 0 0 47 0 0 113 2
238 263
188 263
1 2 2 0 0 0 0 48 49 0 0 2
205 660
205 646
1 0 51 0 0 4096 0 49 0 0 154 2
205 629
205 609
1 1 2 0 0 0 0 50 51 0 0 2
405 603
405 599
2 0 52 0 0 4096 0 51 0 0 145 2
405 581
405 567
1 1 2 0 0 0 0 52 53 0 0 4
239 229
239 232
239 232
239 228
2 0 50 0 0 0 0 53 0 0 111 2
239 210
239 198
2 15 53 0 0 4224 0 20 65 0 0 3
498 174
498 359
404 359
2 14 54 0 0 4224 0 21 65 0 0 4
446 175
447 175
447 349
404 349
2 13 55 0 0 12416 0 22 65 0 0 5
391 175
391 213
436 213
436 339
404 339
2 12 56 0 0 12416 0 23 65 0 0 5
337 174
337 223
426 223
426 329
404 329
2 11 57 0 0 8320 0 24 65 0 0 5
285 173
285 236
416 236
416 319
404 319
1 0 50 0 0 0 0 24 0 0 111 2
276 173
276 198
1 0 50 0 0 0 0 23 0 0 111 2
328 174
328 198
1 0 50 0 0 0 0 22 0 0 111 2
382 175
382 198
1 0 50 0 0 0 0 21 0 0 111 2
437 175
437 198
0 1 50 0 0 4224 0 0 20 113 0 3
188 198
489 198
489 174
31 0 50 0 0 0 0 63 0 0 113 3
154 339
188 339
188 329
32 3 50 0 0 0 0 63 25 0 0 4
154 329
188 329
188 172
187 172
29 2 35 0 0 8320 0 63 25 0 0 3
154 359
178 359
178 172
0 1 2 0 0 0 0 0 25 117 0 2
169 261
169 172
34 0 2 0 0 0 0 63 0 0 117 2
154 309
169 309
33 1 2 0 0 0 0 63 54 0 0 5
154 319
169 319
169 261
147 261
147 269
1 8 2 0 0 0 0 55 65 0 0 3
329 383
329 369
341 369
28 2 58 0 0 4224 0 63 65 0 0 4
154 369
258 369
258 309
341 309
27 3 59 0 0 4224 0 63 65 0 0 4
154 379
269 379
269 319
341 319
26 4 60 0 0 4224 0 63 65 0 0 4
154 389
280 389
280 329
341 329
25 5 61 0 0 4224 0 63 65 0 0 4
154 399
292 399
292 339
341 339
24 6 62 0 0 4224 0 63 65 0 0 4
154 409
303 409
303 349
341 349
7 23 63 0 0 12416 0 65 63 0 0 4
341 359
314 359
314 419
154 419
16 1 42 0 0 8320 0 64 56 0 0 3
672 561
676 561
676 489
1 12 2 0 0 0 0 57 64 0 0 4
640 661
719 661
719 601
672 601
8 1 2 0 0 0 0 64 57 0 0 4
608 631
600 631
600 661
640 661
22 13 64 0 0 4224 0 63 64 0 0 4
154 429
744 429
744 591
672 591
21 14 65 0 0 4224 0 63 64 0 0 4
154 439
722 439
722 581
672 581
20 11 66 0 0 4224 0 63 64 0 0 4
154 449
708 449
708 611
672 611
19 10 67 0 0 4224 0 63 64 0 0 4
154 459
693 459
693 621
672 621
18 5 68 0 0 4224 0 63 64 0 0 4
154 469
543 469
543 601
608 601
17 6 69 0 0 4224 0 63 64 0 0 4
154 479
553 479
553 611
608 611
16 3 70 0 0 4224 0 63 64 0 0 4
154 489
565 489
565 581
608 581
15 2 71 0 0 4224 0 63 64 0 0 4
154 499
577 499
577 571
608 571
8 3 72 0 0 4224 0 63 62 0 0 4
154 569
276 569
276 668
379 668
9 6 73 0 0 8320 0 63 62 0 0 4
154 559
287 559
287 698
379 698
10 5 74 0 0 4224 0 63 62 0 0 4
154 549
299 549
299 688
379 688
12 1 2 0 0 0 0 62 58 0 0 4
443 688
462 688
462 740
365 740
11 11 75 0 0 4224 0 63 62 0 0 4
154 538
509 538
509 698
443 698
12 10 76 0 0 4224 0 63 62 0 0 4
154 529
497 529
497 708
443 708
13 14 77 0 0 4224 0 63 62 0 0 4
154 519
460 519
460 668
443 668
14 13 78 0 0 4224 0 63 62 0 0 4
154 509
472 509
472 678
443 678
7 2 79 0 0 12416 0 63 62 0 0 4
154 579
263 579
263 658
379 658
0 0 52 0 0 8320 0 0 0 146 152 3
339 566
339 567
449 567
2 2 52 0 0 0 0 73 74 0 0 6
312 590
312 566
339 566
339 563
338 563
338 592
0 1 80 0 0 8192 0 0 74 150 0 3
339 708
338 708
338 628
0 1 81 0 0 4096 0 0 73 149 0 2
312 648
312 626
1 2 81 0 0 8320 0 62 2 0 0 4
379 648
312 648
312 816
313 816
7 1 80 0 0 8320 0 62 2 0 0 3
379 708
322 708
322 816
8 1 2 0 0 0 0 62 58 0 0 3
379 718
365 718
365 740
1 16 52 0 0 0 0 59 62 0 0 3
449 566
449 648
443 648
3 0 51 0 0 0 0 63 0 0 154 3
154 619
163 619
163 609
4 1 51 0 0 4224 0 63 60 0 0 2
154 609
225 609
1 0 2 0 0 0 0 63 0 0 156 2
154 639
163 639
2 1 2 0 0 0 0 63 61 0 0 3
154 629
163 629
163 661
77
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 26
696 40 720 184
700 44 716 156
26 Z 
L
I
M
I
T
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
384 55 408 179
388 59 404 155
21 G
L
U
.
D
N
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 7
699 888 763 912
703 892 759 908
7 T HOME1
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 7
601 889 665 913
605 893 661 909
7 T ENC.1
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 8
494 887 566 911
498 891 562 907
8 Z HOME 1
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 7
377 888 441 912
381 892 437 908
7 Z ENC.1
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 9
387 839 411 903
391 843 407 891
9 +
5
V
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 16
276 888 348 932
280 892 344 924
16 X LIN. 
ENCODER
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
713 841 729 865
717 845 725 861
1 +
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
724 841 740 865
728 845 736 861
1 S
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
735 840 751 864
739 844 747 860
1 -
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
512 841 528 865
516 845 524 861
1 +
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
523 841 539 865
527 845 535 861
1 S
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
534 842 550 866
538 846 546 862
1 -
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 9
606 841 630 905
610 845 626 893
9 +
5
V
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
618 841 634 865
622 845 630 861
1 -
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
627 841 643 865
631 845 639 861
1 A
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
638 841 654 865
642 845 650 861
1 B
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
400 841 416 865
404 845 412 861
1 -
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
410 840 426 864
414 844 422 860
1 A
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
421 840 437 864
425 844 433 860
1 B
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
315 839 331 863
319 843 327 859
1 B
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
304 839 320 863
308 843 316 859
1 A
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
295 839 311 863
299 843 307 859
1 -
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 9
283 839 307 903
287 843 303 891
9 +
5
V
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 3
102 630 128 645
106 634 127 645
3 GND
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 3
102 619 128 634
106 623 127 634
3 GND
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 3
108 609 128 624
112 613 127 624
3 +5V
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 3
108 600 128 615
112 604 127 615
3 +5V
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 4
102 589 127 604
106 593 126 604
4 +12V
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 8
83 580 128 595
87 584 127 595
8 LIMIT SW
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 3
105 570 128 585
109 574 127 585
3 XAL
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 4
102 560 128 575
106 564 127 575
4 *XAL
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 3
105 550 128 565
109 554 127 565
3 XBL
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 4
102 540 128 555
106 544 127 555
4 *XBL
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 3
105 529 128 544
109 533 127 544
3 ZA1
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 4
102 520 128 535
106 524 127 535
4 *ZA1
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 3
105 510 128 525
109 514 127 525
3 ZB1
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 4
102 500 128 515
106 504 127 515
4 *ZB1
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 3
105 489 128 504
109 493 127 504
3 ZH1
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 4
102 479 128 494
106 483 127 494
4 *ZH1
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 3
105 470 128 485
109 474 127 485
3 TA1
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 4
102 460 128 475
106 464 127 475
4 *TA1
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 3
105 450 128 465
109 454 127 465
3 TB1
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 4
103 440 129 455
107 444 128 455
4 *TB1
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 3
105 430 128 445
109 434 127 445
3 TH1
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 4
102 420 128 435
106 424 127 435
4 *TH1
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 5
95 410 127 425
99 414 126 425
5 VAC 1
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 6
89 400 128 415
93 404 127 415
6 BLOW 1
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 6
89 390 128 405
93 394 127 405
6 GLU DN
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 5
92 380 128 395
96 384 127 395
5 GLUER
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 7
83 370 128 385
87 374 127 385
7 SPARE 1
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 8
80 360 128 375
84 364 127 375
8 LIGHT ON
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 6
90 349 128 364
94 353 127 364
6 VSEN-1
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 3
102 309 128 324
106 313 127 324
3 GND
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 4
103 329 128 344
107 333 127 344
4 +24V
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 4
103 319 128 334
107 323 127 334
4 +24V
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 8
83 339 128 354
87 343 127 354
8 LIMIT SW
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 3
102 300 128 315
106 304 127 315
3 GND
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
160 133 176 157
164 137 172 153
1 -
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
170 132 186 156
174 136 182 152
1 S
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
180 132 196 156
184 136 192 152
1 +
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 13
266 87 290 171
270 91 286 155
13 +
2
4
V
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
279 55 303 179
283 59 299 155
21 S
P
A
R
E
1
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 13
319 88 343 172
323 92 339 156
13 +
2
4
V
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 17
330 73 354 177
334 77 350 157
17 G
L
U
E
R
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
372 88 396 172
376 92 392 156
13 +
2
4
V
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
428 88 452 172
432 92 448 156
13 +
2
4
V
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 17
441 72 465 176
445 76 461 156
17 B
L
O
W
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
480 87 504 171
484 91 500 155
13 +
2
4
V
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
492 88 516 172
496 92 512 156
13 V
A
C
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
134 115 222 139
138 119 218 135
10 VAC.SENSOR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
553 88 577 172
557 92 573 156
13 +
1
2
V
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
603 90 627 174
607 94 623 158
13 +
1
2
V
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 17
566 72 590 176
570 76 586 156
17 L
I
G
H
T
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
612 57 636 181
616 61 632 157
21 C
A
M
E
R
A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 26
746 43 770 187
750 47 766 159
26 Z 
L
I
M
I
T
2
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
