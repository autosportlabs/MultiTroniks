CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
20 0 30 100 9
20 78 780 559
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
61 C:\PROGRAM FILES\MICROCODE ENGINEERING\CIRCUITMAKER 6\BOM.DAT
0 7
20 78 780 559
144179218 0
0
6 Title:
5 Name:
10 09-17-1998
0
0
23
7 Ground~
168 609 319 0 1 3
0 0
0
0 0 53344 0
0
4 GND8
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8953 0 0
0
0
7 Ground~
168 399 422 0 1 3
0 0
0
0 0 53344 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
4441 0 0
0
0
7 Ground~
168 123 376 0 1 3
0 0
0
0 0 53344 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3618 0 0
0
0
9 Resistor~
219 100 279 0 1 5
0 0
0
0 0 864 90
2 1k
8 0 22 8
2 R5
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612676
82 0 0 0 1 0 0 0
1 R
6153 0 0
0
0
6 Diode~
219 278 327 0 1 5
0 0
0
0 0 832 180
5 DIODE
-18 -18 17 -10
2 D2
-7 -28 7 -20
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 0 0 0 0
1 D
5394 0 0
0
0
7 Ground~
168 173 225 0 1 3
0 0
0
0 0 53344 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7734 0 0
0
0
9 Resistor~
219 128 95 0 1 5
0 0
0
0 0 864 90
2 1k
8 0 22 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612676
82 0 0 0 1 0 0 0
1 R
9914 0 0
0
0
2 +V
167 128 48 0 1 3
0 0
0
0 0 54240 0
2 5V
-7 -22 7 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3747 0 0
0
0
9 Resistor~
219 261 113 0 1 5
0 0
0
0 0 864 90
2 1k
8 0 22 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612720
82 0 0 0 1 0 0 0
1 R
3549 0 0
0
0
9 Resistor~
219 502 136 0 1 5
0 0
0
0 0 864 90
2 1k
8 0 22 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612676
82 0 0 0 1 0 0 0
1 R
7931 0 0
0
0
7 Ground~
168 277 424 0 1 3
0 0
0
0 0 53344 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9325 0 0
0
0
9 Resistor~
219 666 139 0 1 5
0 0
0
0 0 864 90
2 1k
8 0 22 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612720
82 0 0 0 1 0 0 0
1 R
8903 0 0
0
0
2 +V
167 666 74 0 1 3
0 0
0
0 0 54240 0
2 5V
-7 -22 7 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3834 0 0
0
0
7 Ground~
168 602 224 0 1 3
0 0
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3363 0 0
0
0
7 Ground~
168 447 367 0 1 3
0 0
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7668 0 0
0
0
2 +V
167 502 58 0 1 3
0 0
0
0 0 54240 0
3 12V
-10 -22 11 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
4718 0 0
0
0
7 Ground~
168 258 223 0 1 3
0 0
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3874 0 0
0
0
2 +V
167 261 62 0 1 3
0 0
0
0 0 54240 0
3 12V
-10 -22 11 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
6671 0 0
0
0
14 Opto Isolator~
173 194 327 0 1 9
0 0
0
0 0 880 0
7 OPTOISO
-25 -28 24 -20
2 U4
-7 -38 7 -30
0
0
17 %D %1 %2 %3 %4 %S
0
0
4 DIP6
9

0 1 2 5 4 1 2 5 4 -1610612712
88 0 0 0 1 0 0 0
1 U
3789 0 0
0
0
14 Opto Isolator~
173 210 163 0 1 9
0 0
0
0 0 880 512
7 OPTOISO
-26 -28 23 -20
2 U3
-8 -38 6 -30
0
0
17 %D %1 %2 %3 %4 %S
0
0
4 DIP6
9

0 1 2 5 4 1 2 5 4 -1610612720
88 0 0 0 1 0 0 0
1 U
4871 0 0
0
0
14 Opto Isolator~
173 552 187 0 1 9
0 0
0
0 0 880 512
7 OPTOISO
-26 -28 23 -20
2 U1
-8 -38 6 -30
0
0
17 %D %1 %2 %3 %4 %S
0
0
4 DIP6
9

0 1 2 5 4 1 2 5 4 0
88 0 0 0 1 0 0 0
1 U
3750 0 0
0
0
14 Opto Isolator~
173 549 257 0 1 9
0 0
0
0 0 880 0
7 OPTOISO
-25 -28 24 -20
2 U2
-7 -38 7 -30
0
0
17 %D %1 %2 %3 %4 %S
0
0
4 DIP6
9

0 1 2 5 4 1 2 5 4 0
88 0 0 0 1 0 0 0
1 U
8778 0 0
0
0
6 Diode~
219 450 187 0 1 5
0 0
0
0 0 832 0
5 DIODE
-18 -18 17 -10
2 D1
-7 -28 7 -20
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 0 0 0 0
1 D
538 0 0
0
0
35
1 4 0 0 0 0 0 1 22 0 0 3
609 313
609 269
575 269
1 1 0 0 0 0 0 11 2 0 0 4
277 418
277 384
399 384
399 416
1 2 0 0 0 0 0 3 19 0 0 3
123 370
123 339
166 339
2 0 0 0 0 0 0 4 0 0 0 2
100 261
100 239
1 1 0 0 0 0 0 4 19 0 0 3
100 297
100 315
166 315
1 0 0 0 0 0 0 5 0 0 9 3
288 327
311 327
311 339
2 0 0 0 0 0 0 5 0 0 8 3
268 327
250 327
250 315
3 2 0 0 0 0 0 19 22 0 0 4
220 315
502 315
502 269
521 269
4 1 0 0 0 0 0 19 15 0 0 3
220 339
447 339
447 361
1 4 0 0 0 0 0 6 20 0 0 3
173 219
173 175
182 175
0 0 0 0 0 0 0 0 0 12 0 2
128 151
81 151
1 3 0 0 0 0 0 7 20 0 0 3
128 113
128 151
182 151
2 1 0 0 0 0 0 7 8 0 0 2
128 77
128 57
1 1 0 0 0 0 0 20 9 0 0 3
236 151
261 151
261 131
2 1 0 0 0 0 0 9 18 0 0 2
261 95
261 71
1 1 0 0 0 0 0 10 22 0 0 4
502 154
502 244
521 244
521 245
1 2 0 0 0 0 0 16 10 0 0 2
502 67
502 118
0 0 0 0 0 0 0 0 0 21 0 2
666 245
708 245
0 0 0 0 0 0 0 0 0 0 0 2
340 393
340 432
0 0 0 0 0 0 0 0 0 0 0 2
340 347
340 383
3 1 0 0 0 0 0 22 12 0 0 3
575 245
666 245
666 157
1 2 0 0 0 0 0 13 12 0 0 2
666 83
666 121
1 2 0 0 0 0 0 14 21 0 0 3
602 218
602 199
578 199
1 0 0 0 0 0 0 21 0 0 0 3
578 175
619 175
619 59
0 0 0 0 0 0 0 0 0 0 0 2
340 291
340 338
0 0 0 0 0 0 0 0 0 0 0 2
340 240
340 279
0 0 0 0 0 0 0 0 0 0 0 2
340 198
340 229
0 0 0 0 0 0 0 0 0 0 0 2
340 150
340 189
0 0 0 0 0 0 0 0 0 0 0 2
340 118
340 144
0 0 0 0 0 0 0 0 0 0 0 2
340 75
340 111
0 0 0 0 0 0 0 0 0 0 0 2
340 34
340 62
1 0 0 0 0 0 0 23 0 0 34 3
440 187
419 187
419 199
2 0 0 0 0 0 0 23 0 0 35 3
460 187
480 187
480 175
4 1 0 0 0 0 0 21 17 0 0 3
524 199
258 199
258 217
3 2 0 0 0 0 0 21 20 0 0 2
524 175
236 175
11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
347 144 379 168
351 148 375 164
3 J10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
308 145 332 169
312 149 328 165
2 J9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
325 367 341 391
329 371 337 387
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
323 322 339 346
327 326 335 342
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
323 297 339 321
327 301 335 317
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
324 181 340 205
328 185 336 201
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
324 157 340 181
328 161 336 177
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
80 217 128 241
84 221 124 237
5 AVAIL
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
593 36 633 60
597 40 629 56
4 BUSY
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
53 129 93 153
57 133 89 149
4 BUSY
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
693 245 741 269
697 249 737 265
5 AVAIL
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
