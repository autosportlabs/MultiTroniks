CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 40 9
20 78 780 559
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
61 C:\PROGRAM FILES\MICROCODE ENGINEERING\CIRCUITMAKER 6\BOM.DAT
0 7
20 78 780 559
146276370 80
1
76 Title:
        VIDEO EXTENTION CABLE(LVX2)
        P#217018- 
           
51 MULTITRONIKS
ONE FREDERICK ROAD - WARREN, NJ 07059
10 09-17-1998
0
0
2
6 DB-15~
219 854 318 0 15 31
0 2 3 4 5 6 7 8 9 10
11 12 13 14 15 16
0
0 0 2144 512
4 CONN
30 2 58 10
2 J1
-7 -62 7 -54
0
0
0
0
0
6 DB15/F
31

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 1 2 3 4
5 6 7 8 9 10 11 12 13 14
15 0
0 0 0 512 1 1 0 0
1 J
8953 0 0
0
0
3 BNC
94 197 325 0 1 3
0 0
3 BNC
3 0 128 0
0
2 U1
-15 -38 -1 -30
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 0 0 0 0
1 J
4441 0 0
0
0
9
0 0 0 0 0 0 0 0 0 9 7 3
756 322
756 345
817 345
14 0 0 0 0 0 0 1 0 0 7 2
832 300
817 300
13 0 0 0 0 0 0 1 0 0 7 2
832 309
817 309
12 0 0 0 0 0 0 1 0 0 7 2
832 318
817 318
11 0 0 0 0 0 0 1 0 0 7 2
832 327
817 327
10 0 0 0 0 0 0 1 0 0 7 2
832 336
817 336
15 9 0 0 0 0 0 1 1 0 0 4
832 291
817 291
817 345
832 345
0 6 0 0 0 0 0 0 1 9 0 6
782 319
800 319
800 248
884 248
884 304
876 304
0 0 0 0 0 0 0 0 0 0 0 4
234 316
782 316
782 322
233 322
4
-16 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 14
752 383 902 409
756 387 896 405
14 COVER P#17388-
-16 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 29
759 201 959 249
763 205 953 241
29 15 PIN DB CONNECTOR
P#17357-
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 41
355 274 539 318
359 278 535 310
41 CO.AXLE CABLE P#19275-
LENGTH 132 INCHES
-16 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 24
105 231 245 279
109 235 239 271
24 BNC CONNECTOR
P# 17648-
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
