CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
400 190 30 100 9
20 78 780 559
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
61 C:\PROGRAM FILES\MICROCODE ENGINEERING\CIRCUITMAKER 6\BOM.DAT
0 7
20 78 780 559
146276370 80
2
47 Title:SMEEMA INTERFACE CONNECTION (MACHINE END)
50 MULTITRONIKS
ONE FREDERICK ROAD, WARREN, NJ 07059
10 09-17-1998
0
4 LVX2
1
6 CPC14~
94 747 291 0 14 29
0 5 4 3 2 16 17 18 19 20
21 22 23 24 25
6 CPC14~
1 0 4608 0
0
2 U1
73 -5 87 3
0
0
0
0
0
0
29

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 1 2 3 4 5
6 7 8 9 10 11 12 13 14 0
0 0 0 512 1 0 0 0
0
8953 0 0
0
0
14
0 4 2 0 0 4224 0 0 1 0 0 5
181 345
618 345
618 244
703 244
703 264
0 3 3 0 0 4224 0 0 1 0 0 5
182 305
594 305
594 214
778 214
778 240
0 2 4 0 0 4224 0 0 1 0 0 5
183 269
576 269
576 200
747 200
747 240
0 1 5 0 0 4224 0 0 1 0 0 3
182 229
718 229
718 240
0 0 6 0 0 8320 0 0 0 0 0 4
140 200
135 200
135 244
140 244
0 0 7 0 0 8320 0 0 0 0 0 4
140 406
135 406
135 451
140 451
0 0 8 0 0 8320 0 0 0 0 0 4
140 362
135 362
135 285
140 285
0 0 9 0 0 8320 0 0 0 0 0 5
155 406
183 406
183 436
155 436
155 406
0 0 10 0 0 8320 0 0 0 0 0 5
155 368
183 368
183 398
155 398
155 368
0 0 11 0 0 8320 0 0 0 0 0 5
155 330
183 330
183 360
155 360
155 330
0 0 12 0 0 8320 0 0 0 0 0 5
155 292
183 292
183 322
155 322
155 292
0 0 13 0 0 8320 0 0 0 0 0 5
155 254
183 254
183 284
155 284
155 254
0 0 14 0 0 8320 0 0 0 0 0 5
155 215
183 215
183 245
155 245
155 215
0 0 15 0 0 8320 0 0 0 0 0 5
140 200
202 200
202 451
140 451
140 200
8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
703 369 815 393
707 373 811 389
13 CPC 14 FEMALE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 36
114 449 266 493
118 453 262 485
36 HOUSING - 17204-5
TERMINAL - 17205-
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
183 201 199 225
187 205 195 221
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 17
85 171 229 195
89 175 225 191
17 TO CONVEYOR BOARD
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
116 491 292 515
120 495 288 511
21 J9 - TO NEXT CONVEYOR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 26
108 505 324 529
112 509 320 525
26 J10 - TO PREVIOUS CONVEYOR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
344 493 416 517
348 497 412 513
8 LENGTH =
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
344 505 416 529
348 509 412 525
8 LENGTH =
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
