CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
180 280 30 100 9
20 78 780 559
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
61 C:\PROGRAM FILES\MICROCODE ENGINEERING\CIRCUITMAKER 6\BOM.DAT
0 7
20 78 780 559
144179218 80
2
49 Title:SMEEMA INTERFACE CABLE (MACHINE TO MACHINE)
50 MULTITRONIKS
ONE FREDERICK ROAD, WARREN, NJ 07059
10 09-17-1998
0
4 LVX2
2
6 CPC14~
94 721 387 0 14 29
0 5 4 3 2 6 7 8 9 10
11 12 13 14 15
6 CPC14~
1 0 4352 0
5 CPC14
-15 72 20 80
2 U2
73 -5 87 3
0
0
0
0
0
0
29

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 1 2 3 4 5
6 7 8 9 10 11 12 13 14 0
0 0 0 512 1 0 0 0
1 J
8953 0 0
0
0
6 CPC14~
94 257 394 0 14 29
0 5 4 3 2 16 17 18 19 20
21 22 23 24 25
6 CPC14~
2 0 4352 0
6 CPC 14
-19 74 23 82
2 U1
73 -5 87 3
0
0
0
0
0
0
29

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 1 2 3 4 5
6 7 8 9 10 11 12 13 14 0
0 0 0 512 1 0 0 0
1 J
4441 0 0
0
0
4
4 4 2 0 0 8320 0 2 1 0 0 4
213 367
213 265
677 265
677 360
3 3 3 0 0 8320 0 2 1 0 0 4
288 343
288 275
752 275
752 336
2 2 4 0 0 8320 0 2 1 0 0 4
257 343
257 285
721 285
721 336
1 1 5 0 0 8320 0 2 1 0 0 4
228 343
228 296
692 296
692 336
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
749 450 789 474
753 454 785 470
4 MALE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
291 459 331 483
295 463 327 479
4 MALE
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
