CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 10 30 100 9
20 80 780 576
7 5.000 V
7 5.000 V
3 GND
1000 10
24 100 0 1 0
20 Package,Description,
61 C:\PROGRAM FILES\MICROCODE ENGINEERING\CIRCUITMAKER 6\BOM.DAT
0 7
20 80 780 576
143654930 0
0
0
0
0
0
0
48
10 Polar Cap~
219 356 418 0 2 5
0 6 2
0
0 0 832 270
5 2.2uF
12 -1 47 7
2 C5
18 -10 32 -2
0
0
11 %D %1 %2 %V
0
0
7 CapPol1
5

0 1 2 1 2 -1610612559
67 0 0 0 1 0 0 0
1 C
8953 0 0
0
0
7 Ground~
168 284 112 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4441 0 0
0
0
12 NPN Trans:B~
219 387 102 0 3 7
0 2 3 4
0
0 0 832 0
7 MC34064
3 -5 52 3
2 Q5
20 -15 34 -7
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92A
7

0 1 2 3 1 2 3 -1610612676
81 0 0 0 1 0 0 0
1 Q
3618 0 0
0
0
7 Ground~
168 356 443 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6153 0 0
0
0
7 Ground~
168 232 533 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5394 0 0
0
0
7 Ground~
168 168 528 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7734 0 0
0
0
12 NPN Trans:C~
219 177 466 0 3 7
0 11 13 2
0
0 0 832 512
6 2N3904
-64 -1 -22 7
2 Q4
-44 -13 -30 -5
0
0
14 %D %1 %2 %3 %M
0
0
5 TO-39
7

0 1 2 3 1 2 3 -1610612700
81 0 0 0 1 1 0 0
1 Q
9914 0 0
0
0
7 Ground~
168 192 402 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3747 0 0
0
0
7 RSIP10~
219 170 344 0 10 21
0 2 15 16 17 18 22 19 60 20
21
0
0 0 320 90
3 10k
-18 -52 3 -44
3 RN1
-18 -62 3 -54
0
0
125 %DA %1 %2 %V
%DB %1 %3 %V
%DC %1 %4 %V
%DD %1 %5 %V
%DE %1 %6 %V
%DF %1 %7 %V
%DG %1 %8 %V
%DH %1 %9 %V
%DI %1 %10 %V
0
0
5 SIP10
21

0 1 2 3 4 5 6 7 8 9
10 1 2 3 4 5 6 7 8 9
10 -1610612720
82 0 0 512 1 0 0 0
1 R
3549 0 0
0
0
7 Ground~
168 367 180 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7931 0 0
0
0
10 Capacitor~
219 367 154 0 2 5
0 2 3
0
0 0 576 90
15 .01uF CER. CAP.
-30 -5 75 3
2 C2
14 -15 28 -7
0
0
11 %D %1 %2 %V
0
0
7 CapCer1
5

0 1 2 1 2 -1610612704
67 0 0 0 1 0 0 0
1 C
9325 0 0
0
0
7 Ground~
168 487 177 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8903 0 0
0
0
7 Ground~
168 529 168 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3834 0 0
0
0
12 NPN Trans:C~
219 524 105 0 3 7
0 23 26 2
0
0 0 960 0
6 2N3904
22 -2 64 6
2 Q2
36 -12 50 -4
0
0
14 %D %1 %2 %3 %M
0
0
5 TO-39
7

0 1 2 3 1 2 3 -1610612700
81 0 0 0 1 0 0 0
1 Q
3363 0 0
0
0
7 Ground~
168 162 228 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7668 0 0
0
0
10 Capacitor~
219 182 216 0 2 5
0 2 28
0
0 0 576 0
14 18pf CER. CAP.
-50 -18 48 -10
2 C4
-6 10 8 18
0
0
11 %D %1 %2 %V
0
0
7 CapCer1
5

0 1 2 1 2 -1610612676
67 0 0 0 1 0 0 0
1 C
4718 0 0
0
0
10 Capacitor~
219 179 157 0 2 5
0 2 29
0
0 0 576 0
14 18pf CER. CAP.
-49 -18 49 -10
2 C3
-7 -19 7 -11
0
0
11 %D %1 %2 %V
0
0
7 CapCer1
5

0 1 2 1 2 -1610612676
67 0 0 0 1 0 0 0
1 C
3874 0 0
0
0
8 Crystal~
219 207 185 0 2 5
0 28 29
0
0 0 576 90
8 4.000MHZ
13 -5 69 3
3 XL1
-30 -6 -9 2
0
0
11 %D %1 %2 %S
0
32 alias:XCRYSTAL {FREQ=1E6 RS=540}
5 XTAL1
5

0 1 2 1 2 0
88 0 0 0 1 0 0 0
4 XTAL
6671 0 0
0
0
7 Ground~
168 86 329 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3789 0 0
0
0
7 Ground~
168 600 481 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4871 0 0
0
0
7 Ground~
168 434 447 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3750 0 0
0
0
4 LED~
171 504 284 0 2 2
10 30 7
0
0 0 624 0
15 RED LED 5MM/3MM
-76 -4 29 4
2 D1
-24 4 -10 12
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
8778 0 0
0
0
7 Ground~
168 504 442 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
538 0 0
0
0
12 NPN Trans:C~
219 499 368 0 3 7
0 7 25 2
0
0 0 832 0
6 2N3904
14 9 56 17
2 Q1
28 -1 42 7
0
0
14 %D %1 %2 %3 %M
0
0
5 TO-39
7

0 1 2 3 1 2 3 -1610612704
81 0 0 0 1 1 0 0
1 Q
6843 0 0
0
0
7 Ground~
168 74 202 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3136 0 0
0
0
7 Ground~
168 564 244 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5950 0 0
0
0
10 Polar Cap~
219 76 172 0 2 5
0 3 2
0
0 0 576 270
15 10uF ELEC. CAPA
-31 -1 74 7
2 C1
14 -11 28 -3
0
0
11 %D %1 %2 %V
0
0
7 CapPol1
5

0 1 2 1 2 -1610612720
67 0 0 0 1 0 0 0
1 C
5670 0 0
0
0
7 Ground~
168 266 312 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6828 0 0
0
0
4 CON2
94 59 61 0 2 5
0 12 23
4 CON2
1 0 4608 0
15 HEADER 2 PIN MO
-56 -30 49 -22
2 J1
-11 -40 3 -32
0
0
0
0
0
6 MOLEX2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 J
6735 0 0
0
0
4 CON2
94 594 61 0 2 5
0 12 23
4 CON2
2 0 4608 512
15 HEADER 2 PIN MO
-56 -30 49 -22
2 J2
-11 -40 3 -32
0
0
0
0
0
6 MOLEX2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 J
8365 0 0
0
0
4 CON3
94 661 397 0 3 7
0 2 7 8
4 CON3
3 0 4608 0
15 HEADER 3 PIN MO
-48 -31 57 -23
2 J3
-3 -41 11 -33
0
0
0
0
0
6 MOLEX3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 J
4132 0 0
0
0
4 CON3
94 672 288 0 3 7
0 5 10 9
4 CON3
4 0 4608 0
2 TP
-3 -31 11 -23
3 TP1
-6 -41 15 -33
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 J
4551 0 0
0
0
3 REG
94 566 191 0 3 7
0 27 2 3
3 REG
5 0 6912 512
13 5V REG  78L05
-46 -14 45 -6
2 Q3
-5 -24 9 -16
0
0
0
0
0
5 TO-39
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 Q
3635 0 0
0
0
6 VACSEN
94 63 269 0 6 13
0 113 3 5 2 114 115
6 VACSEN
6 0 2560 90
15 PRESSURE SENSOR
-54 -30 51 -22
2 S1
-8 -40 6 -32
0
0
0
0
0
7 VAC SEN
13

0 1 2 3 4 5 6 1 2 3
4 5 6 0
0 0 0 512 1 0 0 0
1 J
3973 0 0
0
0
8 PIC16C71
94 310 239 0 18 37
0 29 28 3 24 2 10 6 9 17
16 15 4 18 22 19 14 20 21
8 PIC16C71
7 0 6272 0
8 PIC16C71
-28 -69 28 -61
2 U1
-7 -79 7 -71
0
0
0
0
0
5 DIP18
37

0 16 15 14 6 5 7 17 8 1
2 3 4 9 10 11 12 13 18 16
15 14 6 5 7 17 8 1 2 3
4 9 10 11 12 13 18 0
0 0 0 0 1 1 0 0
1 U
3851 0 0
0
0
4 CON2
94 75 440 0 2 5
0 11 12
4 CON2
8 0 4736 0
4 CON2
-20 -30 8 -22
2 J4
-13 -40 1 -32
0
0
0
0
0
6 MOLEX2
5

0 1 2 1 2 -1610612720
0 0 0 0 1 0 0 0
1 J
8383 0 0
0
0
9 Resistor~
219 304 396 0 2 5
0 6 5
0
0 0 864 180
3 150
-10 -14 11 -6
3 R12
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612675
82 0 0 0 1 0 0 0
1 R
9334 0 0
0
0
9 Resistor~
219 232 500 0 3 5
0 2 13 -1
0
0 0 864 90
3 47k
5 -5 26 3
3 R10
5 -15 26 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612676
82 0 0 0 1 0 0 0
1 R
7471 0 0
0
0
9 Resistor~
219 232 421 0 2 5
0 13 14
0
0 0 864 90
4 2.2k
8 -6 36 2
3 R11
5 -15 26 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612712
82 0 0 0 1 0 0 0
1 R
3334 0 0
0
0
9 Resistor~
219 415 162 0 2 5
0 4 3
0
0 0 864 90
3 10k
5 -5 26 3
2 R9
8 -15 22 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612720
82 0 0 0 1 0 0 0
1 R
3559 0 0
0
0
9 Resistor~
219 487 138 0 4 5
0 26 2 0 -1
0
0 0 864 270
3 47k
7 0 28 8
2 R7
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612676
82 0 0 0 1 0 0 0
1 R
984 0 0
0
0
9 Resistor~
219 462 105 0 2 5
0 9 26
0
0 0 864 0
4 2.2k
-14 -14 14 -6
2 R6
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612671
82 0 0 0 1 0 0 0
1 R
7557 0 0
0
0
9 Resistor~
219 145 102 0 2 5
0 24 23
0
0 0 864 90
4 750k
8 0 36 8
2 R5
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612720
82 0 0 0 1 0 0 0
1 R
3146 0 0
0
0
9 Resistor~
219 231 178 0 2 5
0 28 29
0
0 0 864 90
3 10M
5 0 26 8
2 R1
7 -10 21 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612676
82 0 0 0 1 0 0 0
1 R
5687 0 0
0
0
9 Resistor~
219 504 223 0 2 5
0 30 3
0
0 0 864 90
3 470
-28 6 -7 14
2 R4
-23 -4 -9 4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612720
82 0 0 0 1 0 0 0
1 R
7939 0 0
0
0
9 Resistor~
219 433 336 0 2 5
0 25 10
0
0 0 864 90
3 10k
5 -5 26 3
2 R2
8 -15 22 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612720
82 0 0 0 1 0 0 0
1 R
3308 0 0
0
0
9 Resistor~
219 434 403 0 4 5
0 25 2 0 -1
0
0 0 864 270
3 47k
7 0 28 8
2 R3
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612676
82 0 0 0 1 0 0 0
1 R
3408 0 0
0
0
9 Resistor~
219 628 351 0 2 5
0 8 27
0
0 0 864 90
7 1K/0.5W
1 -4 50 4
2 R8
8 -15 22 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612676
82 0 0 0 1 0 0 0
1 R
9773 0 0
0
0
67
1 1 2 0 0 8320 0 3 2 0 0 4
392 84
392 74
284 74
284 106
2 0 3 0 0 4096 0 3 0 0 37 3
369 102
310 102
310 131
3 0 4 0 0 4096 0 3 0 0 25 3
392 120
392 189
415 189
0 1 5 0 0 8320 0 0 32 8 0 5
268 396
268 467
580 467
580 277
666 277
2 1 2 0 0 0 0 1 4 0 0 4
355 425
355 424
356 424
356 437
1 0 6 0 0 4096 0 1 0 0 7 2
355 408
355 396
1 7 6 0 0 8320 0 37 35 0 0 4
322 396
404 396
404 206
347 206
3 2 5 0 0 0 0 34 37 0 0 4
70 289
246 289
246 396
286 396
0 2 7 0 0 12416 0 0 31 64 0 4
504 330
570 330
570 396
655 396
1 1 2 0 0 0 0 31 20 0 0 3
655 386
600 386
600 475
1 3 8 0 0 4224 0 48 31 0 0 3
628 369
628 406
655 406
0 3 9 0 0 8320 0 0 32 28 0 5
444 226
444 267
651 267
651 297
666 297
2 0 10 0 0 12416 0 32 0 0 29 4
666 287
568 287
568 257
433 257
1 1 11 0 0 4224 0 36 7 0 0 3
82 430
168 430
168 448
0 2 12 0 0 4096 0 0 36 50 0 3
110 51
110 440
82 440
2 0 13 0 0 4096 0 38 0 0 18 2
232 482
232 468
1 1 2 0 0 0 0 38 5 0 0 2
232 518
232 527
2 1 13 0 0 4224 0 7 39 0 0 5
191 466
232 466
232 468
232 468
232 439
3 1 2 0 0 0 0 7 6 0 0 2
168 484
168 522
16 2 14 0 0 8320 0 35 39 0 0 3
273 256
232 256
232 403
11 2 15 0 0 12416 0 35 9 0 0 4
347 256
395 256
395 378
179 378
10 3 16 0 0 12416 0 35 9 0 0 4
347 246
384 246
384 369
179 369
9 4 17 0 0 12416 0 35 9 0 0 4
347 236
374 236
374 360
179 360
2 0 3 0 0 0 0 40 0 0 61 2
415 144
415 131
12 1 4 0 0 8320 0 35 40 0 0 3
347 266
415 266
415 180
0 1 3 0 0 0 0 0 27 61 0 3
126 131
75 131
75 162
13 5 18 0 0 12416 0 35 9 0 0 4
347 276
365 276
365 351
179 351
8 1 9 0 0 0 0 35 42 0 0 3
347 226
444 226
444 105
6 2 10 0 0 0 0 35 46 0 0 3
347 216
433 216
433 318
15 7 19 0 0 8320 0 35 9 0 0 4
273 245
218 245
218 333
179 333
17 9 20 0 0 4224 0 35 9 0 0 4
273 266
196 266
196 315
179 315
18 10 21 0 0 4224 0 35 9 0 0 4
273 276
187 276
187 306
179 306
1 1 2 0 0 0 0 9 8 0 0 3
179 387
192 387
192 396
14 6 22 0 0 12416 0 35 9 0 0 4
347 286
355 286
355 342
179 342
2 3 3 0 0 0 0 45 33 0 0 5
504 205
504 203
528 203
528 203
527 203
2 0 3 0 0 0 0 11 0 0 61 2
367 145
367 131
3 0 3 0 0 0 0 35 0 0 61 2
310 180
310 131
1 0 23 0 0 4096 0 14 0 0 49 2
529 87
529 61
2 0 23 0 0 0 0 43 0 0 49 2
145 84
145 61
1 4 24 0 0 4224 0 43 35 0 0 5
145 120
145 246
191 246
191 236
273 236
2 1 2 0 0 0 0 47 21 0 0 2
434 421
434 441
0 1 25 0 0 8192 0 0 46 62 0 3
434 369
433 369
433 354
2 1 2 0 0 0 0 41 12 0 0 2
487 156
487 171
1 0 26 0 0 4096 0 41 0 0 47 2
487 120
487 105
1 1 2 0 0 0 0 11 10 0 0 2
367 163
367 174
2 1 2 0 0 0 0 33 26 0 0 2
564 225
564 238
2 2 26 0 0 4224 0 42 14 0 0 2
480 105
506 105
3 1 2 0 0 0 0 14 13 0 0 2
529 123
529 162
2 2 23 0 0 4224 0 29 30 0 0 2
66 61
573 61
1 1 12 0 0 4224 0 29 30 0 0 2
66 51
573 51
1 2 27 0 0 8320 0 33 48 0 0 3
601 202
628 202
628 333
1 0 28 0 0 4096 0 18 0 0 58 2
207 196
207 216
2 0 29 0 0 4096 0 18 0 0 59 2
207 174
207 157
1 2 28 0 0 8320 0 44 35 0 0 3
231 196
231 216
273 216
1 2 29 0 0 8320 0 35 44 0 0 5
273 206
264 206
264 157
231 157
231 160
0 1 2 0 0 0 0 0 15 57 0 2
162 216
162 222
1 1 2 0 0 0 0 17 16 0 0 4
170 157
162 157
162 216
173 216
2 1 28 0 0 0 0 16 44 0 0 3
191 216
231 216
231 196
2 2 29 0 0 0 0 17 44 0 0 3
188 157
231 157
231 160
4 1 2 0 0 0 0 34 19 0 0 3
70 279
86 279
86 323
2 2 3 0 0 12416 0 34 45 0 0 7
70 299
126 299
126 131
460 131
460 203
504 203
504 205
2 1 25 0 0 4224 0 24 47 0 0 3
481 368
434 368
434 385
3 1 2 0 0 0 0 24 23 0 0 2
504 386
504 436
2 1 7 0 0 0 0 22 24 0 0 2
504 294
504 350
1 1 30 0 0 4224 0 45 22 0 0 2
504 241
504 274
5 1 2 0 0 0 0 35 28 0 0 3
273 286
266 286
266 306
2 1 2 0 0 0 0 27 25 0 0 4
75 179
75 193
74 193
74 196
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
