CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
280 90 30 100 9
19 79 772 576
7 5.000 V
7 5.000 V
3 GND
1000 10
24 100 0 1 0
20 Package,Description,
65 C:\PROGRAM FILES\MICROCODE ENGINEERING\CIRCUITMAKER 6 PRO\BOM.DAT
0 7
19 79 772 576
146276370 64
2
21 X-ENC. WIRING DIAGRAM
50 MULTITRONIKS
ONE FREDERICK ROAD, WARREN, NJ 07059
10 10-15-1998
0
4 LVX2
29
10 Connector~
94 595 374 0 2 5
0 2 2
10 Connector~
59 0 96 0
0
0
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
8953 0 0
0
0
10 Connector~
94 595 314 0 2 5
0 5 5
10 Connector~
58 0 96 0
0
0
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
4441 0 0
0
0
10 Connector~
94 595 294 0 2 5
0 6 6
10 Connector~
57 0 96 0
0
0
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
3618 0 0
0
0
10 Connector~
94 595 274 0 2 5
0 7 7
10 Connector~
56 0 96 0
0
0
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
6153 0 0
0
0
10 Connector~
94 595 254 0 2 5
0 8 8
10 Connector~
55 0 96 0
0
0
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
5394 0 0
0
0
10 Connector~
94 595 334 0 2 5
0 4 4
10 Connector~
54 0 96 0
0
0
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
7734 0 0
0
0
10 Connector~
94 595 354 0 2 5
0 3 3
10 Connector~
53 0 96 0
0
0
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
9914 0 0
0
0
10 Connector~
94 595 234 0 2 5
0 9 9
10 Connector~
52 0 96 0
0
0
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
3747 0 0
0
0
10 Connector~
94 595 214 0 2 5
0 10 10
10 Connector~
51 0 96 0
0
0
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
3549 0 0
0
0
10 Connector~
94 225 194 0 2 5
0 10 10
10 Connector~
50 0 96 0
0
0
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
7931 0 0
0
0
10 Connector~
94 225 574 0 2 5
0 2 2
10 Connector~
49 0 96 0
0
0
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
9325 0 0
0
0
10 Connector~
94 225 554 0 2 5
0 3 3
10 Connector~
48 0 96 0
0
0
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
8903 0 0
0
0
10 Connector~
94 225 534 0 2 5
0 4 4
10 Connector~
47 0 96 0
0
0
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
3834 0 0
0
0
10 Connector~
94 225 514 0 2 5
0 5 5
10 Connector~
46 0 96 0
0
0
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
3363 0 0
0
0
10 Connector~
94 225 494 0 2 5
0 6 6
10 Connector~
45 0 96 0
0
0
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
7668 0 0
0
0
10 Connector~
94 225 474 0 2 5
0 7 7
10 Connector~
44 0 96 0
0
0
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
4718 0 0
0
0
10 Connector~
94 225 454 0 2 5
0 8 8
10 Connector~
43 0 96 0
0
0
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
3874 0 0
0
0
10 Connector~
94 225 434 0 2 5
0 17 17
10 Connector~
42 0 96 0
0
0
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
6671 0 0
0
0
10 Connector~
94 225 414 0 2 5
0 16 16
10 Connector~
41 0 96 0
0
0
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
3789 0 0
0
0
10 Connector~
94 225 394 0 2 5
0 15 15
10 Connector~
40 0 96 0
0
0
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
4871 0 0
0
0
10 Connector~
94 225 374 0 2 5
0 14 14
10 Connector~
39 0 96 0
0
0
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
3750 0 0
0
0
10 Connector~
94 225 354 0 2 5
0 13 13
10 Connector~
38 0 96 0
0
0
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
8778 0 0
0
0
10 Connector~
94 225 334 0 2 5
0 12 12
10 Connector~
37 0 96 0
0
0
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
538 0 0
0
0
10 Connector~
94 225 314 0 2 5
0 11 11
10 Connector~
36 0 96 0
0
0
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
6843 0 0
0
0
10 Connector~
94 225 294 0 2 5
0 9 9
10 Connector~
35 0 96 0
0
0
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
3136 0 0
0
0
10 Connector~
94 225 274 0 2 5
0 9 9
10 Connector~
34 0 96 0
0
0
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
5950 0 0
0
0
10 Connector~
94 225 254 0 2 5
0 9 9
10 Connector~
33 0 96 0
0
0
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
5670 0 0
0
0
10 Connector~
94 225 234 0 2 5
0 10 10
10 Connector~
32 0 96 0
0
0
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
6828 0 0
0
0
10 Connector~
94 225 214 0 2 5
0 10 10
10 Connector~
31 0 96 0
0
0
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
6735 0 0
0
0
13
2 1 2 0 0 0 0 11 1 0 0 4
237 574
506 574
506 374
583 374
2 1 3 0 0 0 0 12 7 0 0 4
237 554
486 554
486 354
583 354
2 1 4 0 0 0 0 13 6 0 0 4
237 534
466 534
466 334
583 334
2 1 5 0 0 0 0 14 2 0 0 4
237 514
447 514
447 314
583 314
2 1 6 0 0 0 0 15 3 0 0 4
237 494
425 494
425 294
583 294
2 1 7 0 0 0 0 16 4 0 0 4
237 474
405 474
405 274
583 274
2 1 8 0 0 0 0 17 5 0 0 4
237 454
384 454
384 254
583 254
0 1 9 0 0 0 0 0 8 10 0 4
284 274
326 274
326 234
583 234
0 1 10 0 0 0 0 0 9 12 0 2
284 214
583 214
2 0 9 0 0 0 0 26 0 0 11 2
237 274
285 274
2 2 9 0 0 0 0 27 25 0 0 4
237 254
285 254
285 294
237 294
2 0 10 0 0 0 0 29 0 0 13 2
237 214
285 214
2 2 10 0 0 0 0 10 28 0 0 4
237 194
285 194
285 234
237 234
50
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
242 611 426 635
246 615 422 631
22 X MOTOR ENCODER WIRING
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
195 183 211 207
199 187 207 203
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
195 203 211 227
199 207 207 223
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
195 223 211 247
199 227 207 243
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
194 243 210 267
198 247 206 263
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
195 262 211 286
199 266 207 282
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
194 283 210 307
198 287 206 303
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
194 303 210 327
198 307 206 323
1 7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
194 323 210 347
198 327 206 343
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
194 342 210 366
198 346 206 362
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
187 362 211 386
191 366 207 382
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
188 384 212 408
192 388 208 404
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
188 404 212 428
192 408 208 424
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
187 425 211 449
191 429 207 445
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
186 444 210 468
190 448 206 464
2 14
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
187 462 211 486
191 466 207 482
2 15
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
187 482 211 506
191 486 207 502
2 16
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
186 503 210 527
190 507 206 523
2 17
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
187 522 211 546
191 526 207 542
2 18
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
187 542 211 566
191 546 207 562
2 19
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
186 562 210 586
190 566 206 582
2 20
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 37
196 145 348 189
200 149 344 181
37 2CN TERMINAL ON X 
SERVO(SGDA-04AS)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 39
573 141 749 185
577 145 745 177
39 ENC. OUT FROM X MOTOR
(COLOR OF WIRES)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
523 218 579 242
527 222 575 238
6 ORANGE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
524 237 572 261
528 241 568 257
5 BROWN
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
524 257 572 281
528 261 568 277
5 WHITE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
605 283 645 307
609 287 641 303
4 BLUE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
605 223 637 247
609 227 633 243
3 RED
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
523 317 571 341
527 321 567 337
5 BLACK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
522 337 578 361
526 341 574 357
6 VIOLET
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
605 244 653 268
609 248 649 264
5 GREEN
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
720 224 736 248
724 228 732 244
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
720 242 736 266
724 246 732 262
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
719 260 735 284
723 264 731 280
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
719 283 735 307
723 287 731 303
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
718 302 734 326
722 306 730 322
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
719 322 735 346
723 326 731 342
1 7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
719 342 735 366
723 346 731 362
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
718 360 734 384
722 364 730 380
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
524 297 556 321
528 301 552 317
3 RED
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
606 263 694 287
610 267 690 283
10 GREEN/BLCK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
605 303 693 327
609 307 689 323
10 BLUE/BLACK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
605 322 661 346
609 326 657 342
6 YELLOW
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
605 342 709 366
609 346 705 362
12 YELLOW/BLACK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
605 361 717 385
609 365 713 381
13 ORANGE/SHIELD
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
604 203 644 227
608 207 640 223
4 GRAY
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
720 205 736 229
724 209 732 225
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
525 197 565 221
529 201 561 217
4 GRAY
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
524 276 564 300
528 280 560 296
4 BLUE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
521 357 569 381
525 361 565 377
5 GREEN
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
