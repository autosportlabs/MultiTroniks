CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
210 550 30 100 9
0 66 799 572
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 1
20 Package,Description,
65 C:\PROGRAM FILES\MICROCODE ENGINEERING\CIRCUITMAKER 6 PRO\BOM.DAT
0 7
0 66 799 572
146276370 0
0
6 Title:
5 Name:
0
0
0
44
7 Ground~
168 478 888 0 1 3
0 2
0
0 0 53344 270
0
5 GND21
-17 -28 18 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8953 0 0
0
0
7 Ground~
168 296 375 0 1 3
0 2
0
0 0 53344 0
0
5 GND20
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4441 0 0
0
0
10 Polar Cap~
219 316 354 0 2 5
0 3 2
0
0 0 576 270
6 14046-
0 4 42 12
2 C5
7 -1 21 7
0
0
11 %D %1 %2 %V
0
0
7 RB.2/.4
5

0 1 2 1 2 -1610612604
67 0 0 0 1 0 0 0
1 C
3618 0 0
0
0
10 Polar Cap~
219 273 354 0 2 5
0 4 2
0
0 0 576 270
6 14046-
0 4 42 12
2 C4
14 -6 28 2
0
0
11 %D %1 %2 %V
0
0
7 RB.2/.4
5

0 1 2 1 2 -1610612604
67 0 0 0 1 0 0 0
1 C
6153 0 0
0
0
10 Capacitor~
219 915 244 0 2 5
0 4 2
0
0 0 576 0
6 13521-
-20 -22 22 -14
2 C3
-7 -38 7 -30
0
0
11 %D %1 %2 %V
0
0
6 RAD0.1
5

0 1 2 1 2 -1610612604
67 0 0 0 1 0 0 0
1 C
5394 0 0
0
0
7 Ground~
168 943 243 0 1 3
0 2
0
0 0 53344 90
0
5 GND19
-17 -28 18 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7734 0 0
0
0
7 Ground~
168 1051 817 0 1 3
0 2
0
0 0 53344 0
0
5 GND18
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9914 0 0
0
0
10 Capacitor~
219 1051 785 0 2 5
0 2 3
0
0 0 832 90
5 .01uF
4 0 39 8
2 C2
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.1
5

0 1 2 1 2 -1610612720
67 0 0 0 1 0 0 0
1 C
3747 0 0
0
0
7 Ground~
168 477 845 0 1 3
0 2
0
0 0 53344 0
0
5 GND17
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3549 0 0
0
0
10 Capacitor~
219 477 818 0 2 5
0 2 3
0
0 0 832 90
6 13521-
-57 4 -15 12
2 C1
-36 -6 -22 2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.1
5

0 1 2 1 2 -1610612720
67 0 0 0 1 0 0 0
1 C
7931 0 0
0
0
6 SIP20~
219 820 966 0 20 41
0 2 35 34 90 2 33 32 87 31
30 29 92 93 94 95 96 97 98 99
100
0
0 0 2656 270
7 17463-4
-27 -97 22 -89
3 J15
95 3 116 11
0
0
0
0
0
5 IDC20
41

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 0
0 0 0 512 1 1 0 0
1 J
9325 0 0
0
0
7 Ground~
168 1106 184 0 1 3
0 2
0
0 0 53344 0
0
5 GND16
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8903 0 0
0
0
7 Ground~
168 792 243 0 1 3
0 2
0
0 0 53344 0
0
5 GND15
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3834 0 0
0
0
7 Ground~
168 564 196 0 1 3
0 2
0
0 0 53344 0
0
5 GND14
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3363 0 0
0
0
6 SIP12~
219 1099 148 0 12 25
0 47 46 45 44 43 42 2 48 4
41 40 101
0
0 0 2656 90
8 17419-12
-29 -61 27 -53
3 J14
-15 -50 6 -42
0
0
0
0
0
5 SIP12
25

0 1 2 3 4 5 6 7 8 9
10 11 12 1 2 3 4 5 6 7
8 9 10 11 12 0
0 0 0 512 1 1 0 0
1 J
7668 0 0
0
0
6 SIP12~
219 632 148 0 12 25
0 59 58 57 56 55 54 2 53 4
52 51 102
0
0 0 2656 90
8 17419-12
-29 -61 27 -53
3 J13
-9 -43 12 -35
0
0
0
0
0
5 SIP12
25

0 1 2 3 4 5 6 7 8 9
10 11 12 1 2 3 4 5 6 7
8 9 10 11 12 0
0 0 0 512 1 1 0 0
1 J
4718 0 0
0
0
6 IDC10~
219 621 975 0 10 21
0 2 3 72 71 70 69 103 104 105
106
0
0 0 2656 90
8 17433-1L
-4 -34 52 -26
3 J12
-59 -9 -38 -1
0
0
0
0
0
5 IDC10
21

0 1 2 3 4 5 6 7 8 9
10 1 2 3 4 5 6 7 8 9
10 0
0 0 0 512 1 1 0 0
1 J
3874 0 0
0
0
7 Ground~
168 183 415 0 1 3
0 2
0
0 0 53344 90
0
5 GND13
-17 -28 18 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6671 0 0
0
0
5 DB-37
94 91 598 0 75 75
0 2 3 79 13 11 8 6 38 36
77 107 108 74 18 81 82 83 4 2
2 3 14 12 9 7 39 37 109 110
75 19 80 17 10 78 2 4 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 -1610612428
5 DB-37
1 0 2560 180
6 17680-
-24 -200 18 -192
3 J11
-14 -210 7 -202
0
0
0
0
0
6 DB37/M
75

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 21 22 23 24 25 26 27 29 30
31 32 33 34 35 28 37 36 1 2
3 4 5 6 7 8 9 10 11 12
13 14 15 16 17 18 19 20 21 22
23 24 25 26 27 29 30 31 32 33
34 35 28 37 36 0
0 0 0 512 1 0 0 0
1 J
3789 0 0
0
0
7 Ground~
168 137 793 0 1 3
0 2
0
0 0 53344 0
0
5 GND12
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4871 0 0
0
0
5 SIP26
94 273 972 0 26 53
0 62 63 148 149 64 72 2 2 2
150 151 152 2 153 154 155 2 2 19
18 80 81 17 82 10 83
5 SIP26
2 0 2560 270
7 17463-5
-22 -24 27 -16
3 J10
124 -6 145 2
0
0
0
0
0
5 IDC26
53

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 21 22 23 24 25 26 1 2 3
4 5 6 7 8 9 10 11 12 13
14 15 16 17 18 19 20 21 22 23
24 25 26 0
0 0 0 512 1 0 0 0
1 J
3750 0 0
0
0
5 DB-37
94 394 527 0 75 75
0 2 3 156 157 158 159 85 29 31
27 67 65 60 63 15 160 71 4 2
2 3 161 162 163 84 164 30 68 66
61 62 16 165 64 28 2 4 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 -1610612428
5 DB-37
3 0 2560 180
6 17680-
-24 -200 18 -192
2 J9
-10 -210 4 -202
0
0
0
0
0
6 DB37/M
75

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 21 22 23 24 25 26 27 29 30
31 32 33 34 35 28 37 36 1 2
3 4 5 6 7 8 9 10 11 12
13 14 15 16 17 18 19 20 21 22
23 24 25 26 27 29 30 31 32 33
34 35 28 37 36 0
0 0 0 512 1 0 0 0
1 J
8778 0 0
0
0
6 26LS32
94 558 852 0 16 33
0 85 84 88 203 76 78 77 2 74
75 73 204 89 70 69 3
6 26LS32
4 0 6816 0
6 10463-
-21 -55 21 -47
2 U3
-7 -58 7 -50
0
0
0
0
0
5 DIP16
33

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 1 2 3
4 5 6 7 8 9 10 11 12 13
14 15 16 0
0 0 0 512 1 0 0 0
1 U
538 0 0
0
0
6 IDC50~
219 1318 526 0 101 101
0 205 2 91 2 206 2 90 2 207
2 49 2 208 2 50 2 209 2 73
2 210 2 211 2 212 2 76 2 213
2 214 2 215 2 89 2 216 2 217
2 218 2 88 2 219 2 220 2 221
2 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 -1610612324
0
0 0 6752 0
7 17463-8
-25 -134 24 -126
2 J8
-8 -144 6 -136
0
0
0
0
0
5 IDC50
101

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 21 22 23 24 25 26 27 28 29
30 31 32 33 34 35 36 37 38 39
40 41 42 43 44 45 46 47 48 49
50 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 21 22 23 24 25 26 27 28 29
30 31 32 33 34 35 36 37 38 39
40 41 42 43 44 45 46 47 48 49
50 0
0 0 0 512 1 1 0 0
1 J
6843 0 0
0
0
7 Ground~
168 1352 664 0 1 3
0 2
0
0 0 53344 0
0
5 GND11
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3136 0 0
0
0
7 Ground~
168 1163 663 0 1 3
0 2
0
0 0 53344 0
0
5 GND10
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5950 0 0
0
0
6 IDC50~
219 1129 527 0 101 101
0 222 2 223 2 224 2 225 2 226
2 227 2 228 2 87 2 229 2 230
2 231 2 232 2 233 2 234 2 235
2 236 2 237 2 238 2 239 2 240
2 241 2 86 2 242 2 243 2 244
2 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 -1610612324
0
0 0 6752 0
7 17463-8
-24 -132 25 -124
2 J7
-7 -142 7 -134
0
0
0
0
0
5 IDC50
101

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 21 22 23 24 25 26 27 28 29
30 31 32 33 34 35 36 37 38 39
40 41 42 43 44 45 46 47 48 49
50 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 21 22 23 24 25 26 27 28 29
30 31 32 33 34 35 36 37 38 39
40 41 42 43 44 45 46 47 48 49
50 0
0 0 0 512 1 1 0 0
1 J
5670 0 0
0
0
6 IDC26~
219 939 437 0 26 53
0 32 245 68 67 66 65 61 60 33
246 247 248 249 250 251 252 253 254 255
256 257 258 259 260 261 262
0
0 0 6752 0
7 17463-5
-24 -84 25 -76
2 J6
-7 -73 7 -65
0
0
0
0
0
5 IDC26
53

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 21 22 23 24 25 26 1 2 3
4 5 6 7 8 9 10 11 12 13
14 15 16 17 18 19 20 21 22 23
24 25 26 0
0 0 0 512 1 1 0 0
1 J
6828 0 0
0
0
6 IDC26~
219 755 398 0 26 53
0 54 263 59 58 57 56 52 51 55
264 265 266 267 42 268 47 46 45 44
41 40 43 269 270 271 272
0
0 0 6752 0
7 17463-5
-24 -83 25 -75
2 J5
-7 -93 7 -85
0
0
0
0
0
5 IDC26
53

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 21 22 23 24 25 26 1 2 3
4 5 6 7 8 9 10 11 12 13
14 15 16 17 18 19 20 21 22 23
24 25 26 0
0 0 0 512 1 1 0 0
1 J
6735 0 0
0
0
6 IDC26~
219 752 667 0 26 53
0 34 273 39 38 37 36 274 275 35
276 277 278 279 22 280 26 25 24 23
21 20 5 281 282 283 284
0
0 0 6752 0
7 17463-5
-47 -71 2 -63
2 J4
-30 -81 -16 -73
0
0
0
0
0
5 IDC26
53

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 21 22 23 24 25 26 1 2 3
4 5 6 7 8 9 10 11 12 13
14 15 16 17 18 19 20 21 22 23
24 25 26 0
0 0 0 512 1 1 0 0
1 J
8365 0 0
0
0
6 IDC50~
219 286 204 0 101 101
0 285 2 286 2 19 2 18 2 17
2 16 2 15 2 287 2 14 2 13
2 12 2 11 2 9 2 8 2 7
2 6 2 288 2 289 2 290 2 291
2 292 2 293 2 294 2 10 2 295
2 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 -1610612324
0
0 0 4704 0
7 17463-8
-25 -124 24 -116
2 J3
-8 -134 6 -126
0
0
0
0
0
5 IDC50
101

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 21 22 23 24 25 26 27 28 29
30 31 32 33 34 35 36 37 38 39
40 41 42 43 44 45 46 47 48 49
50 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 21 22 23 24 25 26 27 28 29
30 31 32 33 34 35 36 37 38 39
40 41 42 43 44 45 46 47 48 49
50 0
0 0 0 512 1 1 0 0
1 J
4132 0 0
0
0
4 2003
94 835 196 0 16 33
0 49 296 297 298 299 300 50 2 48
301 302 303 304 305 53 4
4 2003
5 0 4736 0
6 10395-
-22 -56 20 -48
2 U2
-8 -66 6 -58
0
0
0
0
0
5 DIP16
33

0 1 2 3 4 5 6 7 8 16
15 14 13 12 11 10 9 1 2 3
4 5 6 7 8 16 15 14 13 12
11 10 9 0
0 0 0 512 1 0 0 0
1 U
4551 0 0
0
0
6 26LS32
94 971 790 0 16 33
0 27 28 86 306 307 308 309 2 310
311 312 313 314 315 316 3
6 26LS32
6 0 6816 0
6 10463-
-21 -55 21 -47
2 U1
-7 -65 7 -57
0
0
0
0
0
5 DIP16
33

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 1 2 3
4 5 6 7 8 9 10 11 12 13
14 15 16 0
0 0 0 512 1 0 0 0
1 U
3635 0 0
0
0
6 SIP12~
219 1181 967 0 12 25
0 2 91 26 25 24 23 21 20 2
5 2 22
0
0 0 2656 270
8 17419-12
-29 -61 27 -53
2 J2
64 3 78 11
0
0
0
0
0
5 SIP12
25

0 1 2 3 4 5 6 7 8 9
10 11 12 1 2 3 4 5 6 7
8 9 10 11 12 0
0 0 0 0 1 1 0 0
1 J
3973 0 0
0
0
7 Ground~
168 478 343 0 1 3
0 2
0
0 0 53344 90
0
4 GND9
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3851 0 0
0
0
5 SIP4~
219 68 340 0 4 9
0 4 3 79 2
0
0 0 608 512
6 17628-
2 2 44 10
2 J1
-12 -31 2 -23
0
0
0
0
0
8 CON200-4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
1 J
8383 0 0
0
0
7 Ground~
168 111 379 0 1 3
0 2
0
0 0 53344 0
0
4 GND8
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9334 0 0
0
0
7 Ground~
168 429 720 0 1 3
0 2
0
0 0 53344 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7471 0 0
0
0
7 Ground~
168 121 967 0 1 3
0 2
0
0 0 53344 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3334 0 0
0
0
7 Ground~
168 600 1034 0 1 3
0 2
0
0 0 53344 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3559 0 0
0
0
7 Ground~
168 697 967 0 1 3
0 2
0
0 0 53344 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
984 0 0
0
0
7 Ground~
168 918 841 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7557 0 0
0
0
7 Ground~
168 1086 979 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3146 0 0
0
0
7 Ground~
168 357 119 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5687 0 0
0
0
216
1 8 2 0 0 8192 0 1 23 0 0 3
485 889
485 888
525 888
1 0 3 0 0 4096 0 3 0 0 74 2
315 344
315 336
1 0 4 0 0 4096 0 4 0 0 148 2
272 344
272 327
1 2 2 0 0 0 0 2 3 0 0 3
296 369
315 369
315 361
2 1 2 0 0 0 0 4 2 0 0 3
272 361
272 369
296 369
1 0 4 0 0 0 0 5 0 0 101 3
906 244
895 244
895 230
2 1 2 0 0 0 0 5 6 0 0 2
924 244
936 244
2 0 3 0 0 8192 0 8 0 0 57 3
1051 776
1051 763
1018 763
1 1 2 0 0 0 0 7 8 0 0 2
1051 811
1051 794
2 0 3 0 0 8192 0 10 0 0 61 3
477 809
477 791
512 791
1 1 2 0 0 0 0 9 10 0 0 2
477 839
477 827
11 0 2 0 0 0 0 34 0 0 55 2
1143 963
1143 953
22 10 5 0 0 4224 0 30 34 0 0 3
767 703
1152 703
1152 963
0 0 2 0 0 0 0 0 0 15 38 2
321 114
321 104
6 50 2 0 0 8192 0 31 31 0 0 4
301 114
321 114
321 312
302 312
48 0 2 0 0 0 0 31 0 0 15 2
301 303
321 303
46 0 2 0 0 0 0 31 0 0 15 2
301 294
321 294
44 0 2 0 0 0 0 31 0 0 15 2
302 285
321 285
42 0 2 0 0 0 0 31 0 0 15 2
301 276
321 276
40 0 2 0 0 0 0 31 0 0 15 2
301 267
321 267
38 0 2 0 0 0 0 31 0 0 15 2
301 258
321 258
36 0 2 0 0 0 0 31 0 0 15 2
301 249
321 249
34 0 2 0 0 0 0 31 0 0 15 2
301 240
321 240
32 0 2 0 0 0 0 31 0 0 15 2
301 231
321 231
30 0 2 0 0 0 0 31 0 0 15 2
301 222
321 222
28 0 2 0 0 0 0 31 0 0 15 2
301 213
321 213
26 0 2 0 0 0 0 31 0 0 15 2
301 204
321 204
24 0 2 0 0 0 0 31 0 0 15 2
301 195
321 195
22 0 2 0 0 0 0 31 0 0 15 2
301 186
321 186
20 0 2 0 0 0 0 31 0 0 15 2
301 177
321 177
18 0 2 0 0 0 0 31 0 0 15 2
301 168
321 168
16 0 2 0 0 0 0 31 0 0 15 2
301 159
321 159
14 0 2 0 0 0 0 31 0 0 15 2
301 150
321 150
12 0 2 0 0 0 0 31 0 0 15 2
301 141
321 141
10 0 2 0 0 0 0 31 0 0 15 2
301 132
321 132
8 0 2 0 0 0 0 31 0 0 15 2
301 123
321 123
1 0 2 0 0 0 0 44 0 0 38 3
357 113
357 96
321 96
2 4 2 0 0 0 0 31 31 0 0 4
301 96
321 96
321 105
301 105
7 31 6 0 0 8320 0 19 31 0 0 4
114 536
256 536
256 231
266 231
25 29 7 0 0 8320 0 19 31 0 0 4
114 526
248 526
248 222
266 222
6 27 8 0 0 8320 0 19 31 0 0 4
114 516
239 516
239 213
266 213
24 25 9 0 0 8320 0 19 31 0 0 4
114 506
230 506
230 204
266 204
0 47 10 0 0 4224 0 0 31 157 0 3
172 726
172 303
266 303
23 5 11 0 0 8320 0 31 19 0 0 4
266 195
222 195
222 496
114 496
23 21 12 0 0 8320 0 19 31 0 0 4
114 486
213 486
213 186
266 186
19 4 13 0 0 8320 0 31 19 0 0 4
266 177
205 177
205 476
114 476
22 17 14 0 0 8320 0 19 31 0 0 4
114 466
197 466
197 168
266 168
13 15 15 0 0 16512 0 31 22 0 0 8
266 150
188 150
188 389
308 389
308 803
450 803
450 625
417 625
32 11 16 0 0 16512 0 22 31 0 0 8
417 615
442 615
442 794
316 794
316 397
180 397
180 141
266 141
0 9 17 0 0 4224 0 0 31 155 0 3
162 706
162 132
266 132
7 0 18 0 0 8320 0 31 0 0 152 3
266 123
154 123
154 676
0 5 19 0 0 4224 0 0 31 151 0 3
147 666
147 114
266 114
18 0 4 0 0 4096 0 19 0 0 148 4
114 756
140 756
140 745
139 745
9 0 2 0 0 0 0 34 0 0 55 2
1161 963
1161 953
1 1 2 0 0 0 0 43 34 0 0 4
1086 973
1086 953
1233 953
1233 963
1 8 2 0 0 0 0 42 33 0 0 3
918 835
918 826
938 826
0 16 3 0 0 4096 0 0 33 61 0 6
613 800
913 800
913 725
1018 725
1018 763
1004 763
5 0 2 0 0 0 0 11 0 0 59 2
870 962
870 939
1 1 2 0 0 8192 0 41 11 0 0 4
697 961
697 939
906 939
906 962
0 0 3 0 0 4224 0 0 0 61 74 3
519 791
519 308
455 308
16 2 3 0 0 0 0 23 17 0 0 7
591 825
613 825
613 791
512 791
512 948
601 948
601 956
1 1 2 0 0 0 0 40 17 0 0 3
600 1028
601 1028
601 991
17 0 2 0 0 0 0 21 0 0 68 2
244 960
244 942
18 0 2 0 0 0 0 21 0 0 68 2
235 960
235 942
13 0 2 0 0 0 0 21 0 0 68 2
280 960
280 942
9 0 2 0 0 0 0 21 0 0 68 2
316 960
316 942
8 0 2 0 0 0 0 21 0 0 68 2
325 960
325 942
7 1 2 0 0 8192 0 21 39 0 0 4
334 960
334 942
121 942
121 961
0 9 4 0 0 4096 0 0 16 70 0 3
510 299
657 299
657 161
0 0 4 0 0 8320 0 0 0 71 148 5
431 675
510 675
510 299
341 299
341 328
37 18 4 0 0 0 0 22 22 0 0 4
417 675
431 675
431 685
417 685
1 0 2 0 0 0 0 38 0 0 73 2
429 714
429 705
19 36 2 0 0 0 0 22 22 0 0 4
417 705
429 705
429 695
417 695
2 0 3 0 0 0 0 36 0 0 76 8
74 336
349 336
349 337
349 337
349 308
455 308
455 365
435 365
1 4 2 0 0 0 0 37 36 0 0 3
111 373
111 354
74 354
2 21 3 0 0 0 0 22 22 0 0 4
417 365
435 365
435 375
417 375
0 1 2 0 0 0 0 0 35 78 0 3
432 345
432 344
471 344
20 1 2 0 0 0 0 22 22 0 0 4
417 355
432 355
432 345
417 345
21 8 20 0 0 12416 0 30 34 0 0 5
732 703
712 703
712 886
1170 886
1170 963
7 20 21 0 0 8320 0 34 30 0 0 3
1179 963
1179 694
767 694
12 14 22 0 0 8320 0 34 30 0 0 3
1134 963
1134 667
767 667
6 19 23 0 0 8320 0 34 30 0 0 5
1188 963
1188 878
676 878
676 694
732 694
18 5 24 0 0 4224 0 30 34 0 0 3
767 685
1197 685
1197 963
4 17 25 0 0 8320 0 34 30 0 0 5
1206 963
1206 861
684 861
684 685
732 685
3 16 26 0 0 8320 0 34 30 0 0 3
1215 963
1215 676
767 676
10 1 27 0 0 12416 0 22 33 0 0 4
417 525
628 525
628 763
938 763
2 35 28 0 0 4224 0 33 22 0 0 4
938 772
618 772
618 515
417 515
8 11 29 0 0 8320 0 22 11 0 0 3
417 485
816 485
816 962
10 27 30 0 0 8320 0 11 22 0 0 4
825 962
826 962
826 495
417 495
9 9 31 0 0 8320 0 22 11 0 0 3
417 505
834 505
834 962
1 7 32 0 0 16512 0 28 11 0 0 5
919 383
897 383
897 603
852 603
852 962
9 6 33 0 0 16512 0 28 11 0 0 5
919 419
888 419
888 615
861 615
861 962
3 1 34 0 0 8320 0 11 30 0 0 5
888 962
888 789
702 789
702 613
732 613
9 2 35 0 0 12416 0 30 11 0 0 5
732 649
693 649
693 780
897 780
897 962
9 6 36 0 0 12416 0 19 30 0 0 6
114 576
270 576
270 755
797 755
797 631
767 631
27 5 37 0 0 12416 0 19 30 0 0 6
114 566
279 566
279 745
608 745
608 631
732 631
4 8 38 0 0 12416 0 30 19 0 0 6
767 622
807 622
807 736
288 736
288 556
114 556
3 26 39 0 0 12416 0 30 19 0 0 6
732 622
598 622
598 727
299 727
299 546
114 546
11 21 40 0 0 8320 0 15 29 0 0 7
1142 161
1142 282
811 282
811 470
713 470
713 434
735 434
10 20 41 0 0 8320 0 15 29 0 0 5
1133 161
1133 290
820 290
820 425
770 425
0 9 4 0 0 0 0 0 15 111 0 3
873 230
1124 230
1124 161
1 7 2 0 0 0 0 12 15 0 0 2
1106 178
1106 161
14 6 42 0 0 12416 0 29 15 0 0 5
770 398
828 398
828 315
1097 315
1097 161
22 5 43 0 0 12416 0 29 15 0 0 5
770 434
836 434
836 323
1088 323
1088 161
4 19 44 0 0 8320 0 15 29 0 0 5
1079 161
1079 304
706 304
706 425
735 425
3 18 45 0 0 8320 0 15 29 0 0 5
1070 161
1070 332
845 332
845 416
770 416
17 2 46 0 0 12416 0 29 15 0 0 5
735 416
715 416
715 296
1061 296
1061 161
16 1 47 0 0 12416 0 29 15 0 0 5
770 407
854 407
854 341
1052 341
1052 161
9 8 48 0 0 12416 0 32 15 0 0 5
866 160
892 160
892 219
1115 219
1115 161
1 11 49 0 0 12416 0 32 24 0 0 6
803 160
773 160
773 262
1215 262
1215 463
1298 463
0 16 4 0 0 0 0 0 32 69 0 6
657 176
744 176
744 129
873 129
873 230
866 230
1 8 2 0 0 0 0 13 32 0 0 3
792 237
792 230
803 230
15 7 50 0 0 12416 0 24 32 0 0 6
1298 481
1206 481
1206 256
780 256
780 220
803 220
8 11 51 0 0 12416 0 29 16 0 0 5
770 371
794 371
794 267
675 267
675 161
7 10 52 0 0 8320 0 29 16 0 0 3
735 371
666 371
666 161
15 8 53 0 0 12416 0 32 16 0 0 5
866 220
882 220
882 274
648 274
648 161
1 7 2 0 0 0 0 14 16 0 0 4
564 190
564 178
639 178
639 161
1 6 54 0 0 8320 0 29 16 0 0 3
735 344
630 344
630 161
9 5 55 0 0 8320 0 29 16 0 0 3
735 380
621 380
621 161
4 6 56 0 0 8320 0 16 29 0 0 5
612 161
612 281
786 281
786 362
770 362
3 5 57 0 0 4224 0 16 29 0 0 3
603 161
603 362
735 362
4 2 58 0 0 12416 0 29 16 0 0 5
770 353
778 353
778 288
594 288
594 161
1 3 59 0 0 4224 0 16 29 0 0 3
585 161
585 353
735 353
13 8 60 0 0 4224 0 22 28 0 0 4
417 585
981 585
981 410
954 410
30 7 61 0 0 4224 0 22 28 0 0 4
417 575
880 575
880 410
919 410
31 1 62 0 0 8320 0 22 21 0 0 5
417 595
483 595
483 784
388 784
388 959
14 2 63 0 0 16512 0 22 21 0 0 5
417 605
475 605
475 775
379 775
379 960
5 34 64 0 0 4224 0 21 22 0 0 5
352 960
352 764
467 764
467 655
417 655
12 6 65 0 0 4224 0 22 28 0 0 4
417 565
988 565
988 401
954 401
29 5 66 0 0 4224 0 22 28 0 0 4
417 555
872 555
872 401
919 401
11 4 67 0 0 4224 0 22 28 0 0 4
417 545
996 545
996 392
954 392
28 3 68 0 0 4224 0 22 28 0 0 4
417 535
863 535
863 392
919 392
6 15 69 0 0 4224 0 17 23 0 0 3
619 956
619 834
591 834
5 14 70 0 0 12416 0 17 23 0 0 5
619 991
619 999
657 999
657 843
591 843
17 4 71 0 0 8320 0 22 17 0 0 5
417 665
459 665
459 941
610 941
610 956
6 3 72 0 0 16512 0 21 17 0 0 6
343 960
343 952
440 952
440 1000
610 1000
610 991
11 19 73 0 0 4224 0 23 24 0 0 4
591 870
1257 870
1257 499
1298 499
13 9 74 0 0 12416 0 19 23 0 0 6
114 656
234 656
234 934
609 934
609 888
591 888
30 10 75 0 0 12416 0 19 23 0 0 6
114 646
243 646
243 926
601 926
601 879
591 879
27 5 76 0 0 12416 0 24 23 0 0 6
1298 535
1265 535
1265 911
503 911
503 861
525 861
10 7 77 0 0 8320 0 19 23 0 0 4
114 596
252 596
252 879
525 879
35 6 78 0 0 8320 0 19 23 0 0 4
114 586
261 586
261 870
525 870
3 3 79 0 0 8320 0 36 19 0 0 4
74 345
133 345
133 456
114 456
21 0 3 0 0 0 0 19 0 0 147 3
114 446
125 446
125 436
20 0 2 0 0 0 0 19 0 0 146 3
114 426
125 426
125 416
1 1 2 0 0 0 0 19 18 0 0 2
114 416
176 416
0 2 3 0 0 0 0 0 19 74 0 3
349 337
349 436
114 436
1 37 4 0 0 0 0 36 19 0 0 6
74 327
341 327
341 445
139 445
139 746
114 746
19 0 2 0 0 0 0 19 0 0 150 2
114 776
137 776
1 36 2 0 0 0 0 20 19 0 0 3
137 787
137 766
114 766
19 31 19 0 0 0 0 21 19 0 0 3
226 960
226 666
114 666
14 20 18 0 0 0 0 19 21 0 0 3
114 676
217 676
217 960
21 32 80 0 0 4224 0 21 19 0 0 3
208 960
208 686
114 686
15 22 81 0 0 8320 0 19 21 0 0 3
114 696
199 696
199 960
23 33 17 0 0 0 0 21 19 0 0 3
190 960
190 706
114 706
16 24 82 0 0 8320 0 19 21 0 0 3
114 716
181 716
181 960
25 34 10 0 0 0 0 21 19 0 0 3
172 960
172 726
114 726
26 17 83 0 0 4224 0 21 19 0 0 3
163 960
163 736
114 736
2 25 84 0 0 8320 0 23 22 0 0 4
525 834
492 834
492 455
417 455
7 1 85 0 0 8320 0 22 23 0 0 4
417 465
501 465
501 825
525 825
43 3 86 0 0 4224 0 27 33 0 0 4
1109 608
925 608
925 781
938 781
15 8 87 0 0 16512 0 27 11 0 0 5
1109 482
973 482
973 593
843 593
843 962
0 2 2 0 0 0 0 0 27 165 0 3
1163 428
1163 419
1144 419
6 0 2 0 0 0 0 27 0 0 165 2
1144 437
1163 437
4 1 2 0 0 8192 0 27 26 0 0 3
1144 428
1163 428
1163 657
50 0 2 0 0 0 0 27 0 0 165 2
1145 635
1163 635
48 0 2 0 0 0 0 27 0 0 165 2
1144 626
1163 626
46 0 2 0 0 0 0 27 0 0 165 2
1144 617
1163 617
44 0 2 0 0 0 0 27 0 0 165 2
1145 608
1163 608
42 0 2 0 0 0 0 27 0 0 165 2
1144 599
1163 599
40 0 2 0 0 0 0 27 0 0 165 2
1144 590
1163 590
38 0 2 0 0 0 0 27 0 0 165 2
1144 581
1163 581
36 0 2 0 0 0 0 27 0 0 165 2
1144 572
1163 572
34 0 2 0 0 0 0 27 0 0 165 2
1144 563
1163 563
32 0 2 0 0 0 0 27 0 0 165 2
1144 554
1163 554
30 0 2 0 0 0 0 27 0 0 165 2
1144 545
1163 545
28 0 2 0 0 0 0 27 0 0 165 2
1144 536
1163 536
26 0 2 0 0 0 0 27 0 0 165 2
1144 527
1163 527
24 0 2 0 0 0 0 27 0 0 165 2
1144 518
1163 518
22 0 2 0 0 0 0 27 0 0 165 2
1144 509
1163 509
20 0 2 0 0 0 0 27 0 0 165 2
1144 500
1163 500
18 0 2 0 0 0 0 27 0 0 165 2
1144 491
1163 491
16 0 2 0 0 0 0 27 0 0 165 2
1144 482
1163 482
14 0 2 0 0 0 0 27 0 0 165 2
1144 473
1163 473
12 0 2 0 0 0 0 27 0 0 165 2
1144 464
1163 464
10 0 2 0 0 0 0 27 0 0 165 2
1144 455
1163 455
8 0 2 0 0 0 0 27 0 0 165 2
1144 446
1163 446
43 3 88 0 0 12416 0 24 23 0 0 6
1298 607
1272 607
1272 918
492 918
492 843
525 843
35 13 89 0 0 12416 0 24 23 0 0 4
1298 571
1248 571
1248 852
591 852
7 4 90 0 0 12416 0 24 11 0 0 5
1298 445
1231 445
1231 648
879 648
879 962
3 2 91 0 0 8320 0 24 34 0 0 3
1298 427
1224 427
1224 963
0 2 2 0 0 0 0 0 24 194 0 3
1352 427
1352 418
1333 418
6 0 2 0 0 0 0 24 0 0 194 2
1333 436
1352 436
4 1 2 0 0 8320 0 24 25 0 0 3
1333 427
1352 427
1352 658
50 0 2 0 0 0 0 24 0 0 194 2
1334 634
1352 634
48 0 2 0 0 0 0 24 0 0 194 2
1333 625
1352 625
46 0 2 0 0 0 0 24 0 0 194 2
1333 616
1352 616
44 0 2 0 0 0 0 24 0 0 194 2
1334 607
1352 607
42 0 2 0 0 0 0 24 0 0 194 2
1333 598
1352 598
40 0 2 0 0 0 0 24 0 0 194 2
1333 589
1352 589
38 0 2 0 0 0 0 24 0 0 194 2
1333 580
1352 580
36 0 2 0 0 0 0 24 0 0 194 2
1333 571
1352 571
34 0 2 0 0 0 0 24 0 0 194 2
1333 562
1352 562
32 0 2 0 0 0 0 24 0 0 194 2
1333 553
1352 553
30 0 2 0 0 0 0 24 0 0 194 2
1333 544
1352 544
28 0 2 0 0 0 0 24 0 0 194 2
1333 535
1352 535
26 0 2 0 0 0 0 24 0 0 194 2
1333 526
1352 526
24 0 2 0 0 0 0 24 0 0 194 2
1333 517
1352 517
22 0 2 0 0 0 0 24 0 0 194 2
1333 508
1352 508
20 0 2 0 0 0 0 24 0 0 194 2
1333 499
1352 499
18 0 2 0 0 0 0 24 0 0 194 2
1333 490
1352 490
16 0 2 0 0 0 0 24 0 0 194 2
1333 481
1352 481
14 0 2 0 0 0 0 24 0 0 194 2
1333 472
1352 472
12 0 2 0 0 0 0 24 0 0 194 2
1333 463
1352 463
10 0 2 0 0 0 0 24 0 0 194 2
1333 454
1352 454
8 0 2 0 0 0 0 24 0 0 194 2
1333 445
1352 445
70
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
29 344 57 364
33 348 54 362
3 GND
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 4
22 336 57 356
26 340 54 354
4 +12V
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
28 326 56 346
32 330 53 344
3 +5V
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 4
22 316 57 336
26 320 54 334
4 +24V
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 310
734 998 914 1209
738 1001 911 1170
310 PIN             DES
-------------------------
1               GND
2               Z REF(+)
3               Z REF(-)
4               Z INH
5               GND
6               B REF(+)
7               B REF(-)
8               B INH
9               HALL 1
10              HALL 2
11              HALL 3
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 280
282 982 443 1240
286 986 440 1196
280 PIN         DES
--------------------
14          
15         
16          
17          GND 
18          GND
19          VAC 1
20          BLOW 1
21          GLU DWN
22          GLU ON
23          SPARE 1
24          LIGHT ON
25          VAC SEN 1
26          LIMIT 1
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 265
118 982 265 1240
122 986 262 1196
265 PIN         DES
-----------------
1           VAC 2
2           BLOW 2
3           SPARE 2
4           SPARE 3
5           V SEN 2
6           LIMIT 2
7           GND
8           GND
9           GND
10         
11          
12         
13          GND
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 222
1125 1002 1300 1243
1129 1006 1297 1202
222 PIN            DES
-----------------------
1          EN GND
2          EN +
3          A+
4          A-
5          B+
6          B-
7          IND+
8          IND-
9
10
11         +/-ANALOG
12         ANA.GND
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
1165 980 1207 1000
1169 984 1204 998
5 THETA
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
328 573 370 593
332 577 367 591
5 *BIND
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 4
335 564 370 584
339 568 367 582
4 BIND
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 4
335 583 370 603
339 587 367 601
4 VAC2
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
328 594 370 614
332 598 367 612
5 BLOW2
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
328 643 370 663
332 647 367 661
5 VSEN2
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 4
334 655 369 675
338 659 366 673
4 L SW
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
342 556 370 576
346 560 367 574
3 *BB
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
349 545 370 565
353 549 367 563
2 BB
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
342 534 370 554
346 538 367 552
3 *BA
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
348 523 369 543
352 527 366 541
2 BA
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
329 444 369 463
333 447 366 460
5 XHOME
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
322 454 369 473
326 457 366 470
6 *XHOME
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
314 492 370 516
318 496 366 512
6 HALL 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
314 471 370 495
318 475 366 491
6 HALL 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
314 481 370 505
318 485 366 501
6 HALL 2
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
328 504 370 524
332 508 367 522
5 BHOME
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
321 514 370 534
325 518 367 532
6 *BHOME
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
1072 105 1121 125
1076 109 1118 123
6 Y AXIS
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
608 111 657 131
612 115 654 129
6 X AXIS
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 11
575 1001 659 1021
579 1005 656 1019
11 Y INTERFACE
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 4
1259 469 1294 489
1263 472 1291 486
4 X EN
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 4
1259 450 1294 470
1263 454 1291 468
4 Y EN
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 4
1260 432 1295 452
1264 436 1292 450
4 Z EN
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 4
1260 414 1295 434
1264 418 1292 432
4 T EN
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
1239 594 1288 614
1243 598 1285 612
6 X HOME
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
1238 558 1287 578
1242 562 1284 576
6 Y HOME
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
1237 522 1286 542
1241 526 1283 540
6 Z HOME
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
1235 486 1284 506
1239 490 1281 504
6 T HOME
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
1051 592 1100 612
1055 596 1097 610
6 B HOME
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 4
1067 469 1102 489
1071 473 1099 487
4 B EN
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
738 457 766 477
742 461 763 475
3 X,Y
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
736 727 764 747
740 731 761 745
3 Z,T
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
929 495 943 515
933 499 940 513
1 B
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
47 537 68 557
51 541 65 555
2 ZA
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
40 546 68 566
44 550 65 564
3 *ZA
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
47 556 68 576
51 560 65 574
2 ZB
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
40 566 68 586
44 570 65 584
3 *ZB
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
26 576 68 596
30 580 65 594
5 ZHOME
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
19 585 68 605
23 589 65 603
6 *ZHOME
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
46 595 67 615
50 599 64 613
2 TA
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
40 604 68 624
44 608 65 622
3 *TA
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
47 615 68 635
51 619 65 633
2 TB
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
40 625 68 645
44 629 65 643
3 *TB
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
27 634 69 654
31 638 66 652
5 THOME
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
20 643 69 663
24 647 66 661
6 *THOME
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 4
34 654 69 674
38 658 66 672
4 VAC1
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
28 664 70 684
32 668 67 682
5 BLOW1
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
27 674 69 694
31 678 66 692
5 GLUDN
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
27 684 69 704
31 688 66 702
5 GLUER
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
21 695 70 715
25 699 67 713
6 SPARE1
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 7
14 705 70 725
18 709 67 723
7 LIGHTON
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
28 715 70 735
32 719 67 733
5 VSEN1
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
28 725 70 745
32 729 67 743
5 LIMIT
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
704 330 732 350
708 334 729 348
3 GND
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 10
665 365 742 385
669 369 739 383
10 +/-10V AN.
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
651 366 665 386
655 370 662 384
1 X
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
771 383 799 403
775 387 796 401
3 GND
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 10
963 311 1040 331
967 315 1037 329
10 +/-10V AN.
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
952 312 966 332
956 316 963 330
1 Y
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 4
825 977 856 1000
830 982 855 997
4 BETA
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
883 977 895 1000
888 982 894 997
1 Z
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
