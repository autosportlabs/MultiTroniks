CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 40 9
20 78 780 559
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
61 C:\PROGRAM FILES\MICROCODE ENGINEERING\CIRCUITMAKER 6\BOM.DAT
0 7
20 78 780 559
146276370 80
2
25 Title:VIDEO MONITOR CABLE
56 Name:MULTITRONIKS
ONE FREDERICK ROAD - WARREN, NJ 07059
10 09-17-1998
0
0
2
3 BNC
94 850 388 0 1 3
0 0
3 BNC
5 0 128 512
0
2 U2
-15 -38 -1 -30
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 0 0 0 0
1 J
8953 0 0
0
0
3 BNC
94 147 388 0 1 3
0 0
3 BNC
4 0 128 0
0
2 U1
-15 -38 -1 -30
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 0 0 0 0
1 J
4441 0 0
0
0
2
0 0 0 0 0 0 0 0 0 0 0 2
183 386
798 386
0 0 0 0 0 0 0 0 0 0 0 2
183 380
799 380
3
-16 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 23
81 316 221 364
85 320 215 356
23 BNC CONNECTOR
P#17648-
-16 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 23
799 318 939 366
803 322 933 358
23 BNC CONNECTOR
P#17648-
-16 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 41
285 339 525 387
289 343 519 379
41 CO.AXLE CABLE P# 19275-
LENGTH 48 INCHES
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
