CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 15 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 10 10 13 
10 18 11 
0 10 30 40 9
24 84 784 576
7 5.000 V
7 5.000 V
3 GND
1000 10
24 100 1 1 0
20 Package,Description,
65 C:\PROGRAM FILES\MICROCODE ENGINEERING\CIRCUITMAKER 6 PRO\BOM.DAT
0 7
24 84 784 576
146276370 80
2
20 CONVEYOR ELE. WIRING
51 MULTITRONIKS
ONE FREDERICK ROAD, WARREN, NJ. 07059
10 03-19-1999
1 1
6 LVX II
54
7 ACMOTOR
94 911 332 0 4 9
0 18 17 18 16
7 ACMOTOR
1 0 128 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
0
8953 0 0
0
0
10 Connector~
94 734 304 0 2 5
0 18 18
10 Connector~
2 0 96 180
0
0
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
4441 0 0
0
0
10 Connector~
94 734 317 0 2 5
0 17 17
10 Connector~
3 0 96 180
0
0
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
3618 0 0
0
0
10 Connector~
94 734 329 0 2 5
0 18 18
10 Connector~
4 0 96 180
0
0
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
6153 0 0
0
0
10 Connector~
94 734 341 0 2 5
0 16 16
10 Connector~
5 0 96 180
0
0
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
5394 0 0
0
0
10 Connector~
94 734 354 0 2 5
0 32 32
10 Connector~
6 0 96 180
0
0
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
7734 0 0
0
0
10 Connector~
94 735 367 0 2 5
0 33 33
10 Connector~
7 0 96 180
0
0
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
9914 0 0
0
0
7 ACMOTOR
94 911 435 0 4 9
0 15 14 15 13
7 ACMOTOR
8 0 128 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
0
3747 0 0
0
0
10 Connector~
94 736 407 0 2 5
0 15 15
10 Connector~
9 0 96 180
0
0
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
3549 0 0
0
0
10 Connector~
94 736 420 0 2 5
0 14 14
10 Connector~
10 0 96 180
0
0
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
7931 0 0
0
0
10 Connector~
94 736 432 0 2 5
0 15 15
10 Connector~
11 0 96 180
0
0
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
9325 0 0
0
0
6 Input~
177 545 451 0 17 19
0 2 0 0 0 0 0 0 0 0
65 67 32 49 49 48 86 32
0
0 0 53344 512
0
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8903 0 0
0
0
6 Input~
177 545 431 0 17 19
0 3 0 0 0 0 0 0 0 0
78 101 117 116 114 97 108 32
0
0 0 53344 512
0
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3834 0 0
0
0
10 Capacitor~
219 434 411 0 2 5
0 8 19
0
0 0 320 0
3 2uF
-11 -18 10 -10
2 C1
-8 -28 6 -20
0
0
11 %D %1 %2 %V
0
0
6 CAP0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3363 0 0
0
0
10 Capacitor~
219 433 381 0 2 5
0 10 20
0
0 0 320 0
3 2uF
-11 -18 10 -10
2 C2
-8 -28 6 -20
0
0
11 %D %1 %2 %V
0
0
6 CAP0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7668 0 0
0
0
10 TER BLOCK~
94 480 372 0 2 5
0 10 17
10 TER BLOCK~
12 0 0 0
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 0 1 0 0 0
0
4718 0 0
0
0
10 TER BLOCK~
94 480 382 0 2 5
0 20 16
10 TER BLOCK~
13 0 0 0
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 0 1 0 0 0
0
3874 0 0
0
0
10 TER BLOCK~
94 480 392 0 2 5
0 21 18
10 TER BLOCK~
14 0 0 0
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 0 1 0 0 0
0
6671 0 0
0
0
10 TER BLOCK~
94 480 402 0 2 5
0 8 14
10 TER BLOCK~
15 0 0 0
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 0 1 0 0 0
0
3789 0 0
0
0
10 TER BLOCK~
94 480 412 0 2 5
0 19 13
10 TER BLOCK~
16 0 0 0
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 0 1 0 0 0
0
4871 0 0
0
0
10 TER BLOCK~
94 480 422 0 2 5
0 21 15
10 TER BLOCK~
17 0 0 0
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 0 1 0 0 0
0
3750 0 0
0
0
10 TER BLOCK~
94 480 432 0 2 5
0 21 3
10 TER BLOCK~
18 0 0 0
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 0 1 0 0 0
0
8778 0 0
0
0
10 TER BLOCK~
94 480 442 0 2 5
0 9 2
10 TER BLOCK~
19 0 0 0
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 0 1 0 0 0
0
538 0 0
0
0
10 TER BLOCK~
94 480 452 0 2 5
0 7 2
10 TER BLOCK~
20 0 0 0
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 0 1 0 0 0
0
6843 0 0
0
0
10 Connector~
94 736 444 0 2 5
0 13 13
10 Connector~
21 0 96 180
0
0
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
3136 0 0
0
0
10 Connector~
94 737 458 0 2 5
0 34 34
10 Connector~
22 0 96 180
0
0
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
5950 0 0
0
0
10 Connector~
94 737 472 0 2 5
0 35 35
10 Connector~
23 0 96 180
0
0
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
5670 0 0
0
0
8 Stepper~
185 932 135 0 6 17
13 26 38 25 23 39 24
0
0 0 4192 0
4 100H
10 -16 38 -8
2 L3
17 -26 31 -18
0
0
130 %DA %1 N%DA %V
R%DA N%DA %2 10
%DB %3 N%DB %V
R%DB N%DB %2 10
%DC %4 N%DC %V
R%DC N%DC %5 10
%DD %6 N%DD %V
R%DD N%DD %5 10
0
0
4 SIP6
13

0 1 2 3 4 5 6 1 2 3
4 5 6 0
76 0 0 512 1 0 0 0
1 M
6828 0 0
0
0
10 Connector~
94 753 105 0 2 5
0 26 26
10 Connector~
24 0 96 180
0
0
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
6735 0 0
0
0
7 Output~
178 445 715 0 17 19
0 4 0 0 0 0 0 0 0 0
83 111 108 101 110 111 105 100
0
0 0 53344 0
0
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8365 0 0
0
0
7 Output~
178 445 695 0 17 19
0 4 0 0 0 0 0 0 0 0
83 111 108 101 110 111 105 100
0
0 0 53344 0
0
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4132 0 0
0
0
5 SIP2~
219 324 633 0 2 5
0 4 4
0
0 0 96 90
4 CONN
9 2 37 10
0
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 -1610612616
0 0 0 0 1 0 0 0
1 J
4551 0 0
0
0
5 Ter2~
94 343 497 0 2 5
0 8 7
4 Ter2
25 0 0 0
0
0
0
0
0
0
0
0
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
0
3635 0 0
0
0
5 Ter2~
94 344 377 0 2 5
0 10 9
4 Ter2
26 0 0 0
0
0
0
0
0
0
0
0
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
0
3973 0 0
0
0
6 Input~
177 679 207 0 17 19
0 5 0 0 0 0 0 0 0 0
50 52 86 32 68 67 32 32
0
0 0 53344 512
0
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3851 0 0
0
0
6 Input~
177 679 190 0 17 19
0 6 0 0 0 0 0 0 0 0
48 86 32 32 32 32 32 32
0
0 0 53344 512
0
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8383 0 0
0
0
5 Ter2~
94 594 116 0 2 5
0 26 25
4 Ter2
27 0 0 0
0
0
0
0
0
0
0
0
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
0
9334 0 0
0
0
5 Ter2~
94 594 136 0 2 5
0 23 24
4 Ter2
28 0 0 0
0
0
0
0
0
0
0
0
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
0
7471 0 0
0
0
5 Ter2~
94 594 156 0 2 5
0 6 5
4 Ter2
29 0 0 0
0
0
0
0
0
0
0
0
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
0
3334 0 0
0
0
5 Ter2~
94 491 124 0 2 5
0 30 29
4 Ter2
30 0 0 180
0
0
0
0
0
0
0
0
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
0
3559 0 0
0
0
5 Ter2~
94 491 144 0 2 5
0 40 28
4 Ter2
31 0 0 180
0
0
0
0
0
0
0
0
5

0 1 2 1 2 0
0 0 0 512 1 0 0 0
0
984 0 0
0
0
5 Ter1~
94 157 306 0 1 3
0 30
4 Ter1
32 0 0 90
0
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
7557 0 0
0
0
5 Ter1~
94 167 306 0 1 3
0 29
4 Ter1
33 0 0 90
0
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3146 0 0
0
0
5 Ter1~
94 177 306 0 1 3
0 28
4 Ter1
34 0 0 90
0
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
5687 0 0
0
0
5 SIP 3
94 245 632 0 3 7
0 41 42 43
5 SIP 3
35 0 0 90
4 CONN
-14 -27 14 -19
0
0
0
0
0
0
0
7

0 1 2 3 1 2 3 0
0 0 0 512 1 0 0 0
1 A
7939 0 0
0
0
5 SIP 3
94 189 632 0 3 7
0 44 45 46
5 SIP 3
36 0 0 90
4 CONN
-14 -27 14 -19
0
0
0
0
0
0
0
7

0 1 2 3 1 2 3 0
0 0 0 512 1 0 0 0
1 A
3308 0 0
0
0
5 SIP 3
94 136 632 0 3 7
0 47 48 49
5 SIP 3
37 0 0 90
4 CONN
-14 -27 14 -19
0
0
0
0
0
0
0
7

0 1 2 3 1 2 3 0
0 0 0 512 1 0 0 0
1 A
3408 0 0
0
0
5 SIP 3
94 82 632 0 3 7
0 50 51 52
5 SIP 3
38 0 0 90
4 CONN
-14 -27 14 -19
0
0
0
0
0
0
0
7

0 1 2 3 1 2 3 0
0 0 0 512 1 0 0 0
1 A
9773 0 0
0
0
5 SIP 3
94 33 632 0 3 7
0 53 54 55
5 SIP 3
39 0 0 90
4 CONN
-14 -27 14 -19
0
0
0
0
0
0
0
7

0 1 2 3 1 2 3 0
0 0 0 512 1 0 0 0
1 A
691 0 0
0
0
10 Connector~
94 753 117 0 2 5
0 25 25
10 Connector~
40 0 96 180
0
0
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
7834 0 0
0
0
10 Connector~
94 753 129 0 2 5
0 36 36
10 Connector~
41 0 96 180
0
0
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
3588 0 0
0
0
10 Connector~
94 753 141 0 2 5
0 37 37
10 Connector~
42 0 96 180
0
0
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
4528 0 0
0
0
10 Connector~
94 753 153 0 2 5
0 23 23
10 Connector~
43 0 96 180
0
0
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
3303 0 0
0
0
10 Connector~
94 753 165 0 2 5
0 24 24
10 Connector~
44 0 96 180
0
0
0
0
0
0
0
0
5

0 0 0 0 0 0
0 0 0 0 1 0 0 0
0
9654 0 0
0
0
49
2 1 7 0 0 4224 0 33 24 0 0 4
356 501
420 501
420 451
462 451
1 0 8 0 0 8320 0 33 0 0 24 3
356 491
410 491
410 411
2 1 9 0 0 12416 0 34 23 0 0 4
357 381
400 381
400 441
462 441
0 1 10 0 0 4224 0 0 16 25 0 2
409 371
462 371
0 0 11 0 0 8320 0 0 0 0 0 5
720 393
751 393
751 480
720 480
720 393
0 0 12 0 0 8320 0 0 0 0 0 5
717 282
749 282
749 376
717 376
717 282
2 2 13 0 0 4224 0 25 20 0 0 4
724 444
593 444
593 411
495 411
2 2 14 0 0 4096 0 19 10 0 0 4
495 401
621 401
621 420
724 420
0 2 15 0 0 12288 0 0 11 10 0 4
606 421
607 421
607 432
724 432
2 2 15 0 0 12288 0 21 9 0 0 4
495 421
606 421
606 407
724 407
2 2 16 0 0 4096 0 17 5 0 0 4
495 381
620 381
620 341
722 341
2 2 17 0 0 4096 0 3 16 0 0 4
722 317
598 317
598 371
495 371
2 0 18 0 0 4096 0 4 0 0 14 2
722 329
642 329
2 2 18 0 0 4224 0 18 2 0 0 4
495 391
642 391
642 304
722 304
1 4 13 0 0 0 0 25 8 0 0 2
748 444
875 444
3 1 15 0 0 0 0 8 11 0 0 4
875 430
860 430
860 432
748 432
1 2 14 0 0 4224 0 10 8 0 0 2
748 420
875 420
1 1 15 0 0 4224 0 8 9 0 0 2
875 407
748 407
1 4 16 0 0 4224 0 5 1 0 0 2
746 341
875 341
1 3 18 0 0 0 0 4 1 0 0 4
746 329
860 329
860 327
875 327
1 2 17 0 0 4224 0 3 1 0 0 2
746 317
875 317
1 1 18 0 0 0 0 2 1 0 0 2
746 304
875 304
2 1 19 0 0 4224 0 14 20 0 0 2
443 411
462 411
1 1 8 0 0 0 0 19 14 0 0 4
462 401
410 401
410 411
425 411
1 1 10 0 0 0 0 15 34 0 0 4
424 381
409 381
409 371
357 371
1 2 20 0 0 4224 0 17 15 0 0 2
462 381
442 381
1 0 21 0 0 8320 0 18 0 0 28 3
462 391
449 391
449 421
1 1 21 0 0 0 0 22 21 0 0 4
462 431
449 431
449 421
462 421
2 1 2 0 0 4224 0 24 12 0 0 2
495 451
511 451
2 1 3 0 0 4224 0 22 13 0 0 2
495 431
511 431
2 2 2 0 0 0 0 23 24 0 0 2
495 441
495 451
0 0 22 0 0 8320 0 0 0 0 0 5
737 87
769 87
769 179
737 179
737 87
1 2 23 0 0 12288 0 38 53 0 0 4
607 130
662 130
662 153
741 153
2 2 24 0 0 12288 0 38 54 0 0 4
607 140
648 140
648 165
741 165
1 6 24 0 0 4224 0 54 28 0 0 2
765 165
896 165
1 4 23 0 0 4224 0 53 28 0 0 2
765 153
896 153
2 2 25 0 0 8320 0 37 50 0 0 3
607 120
607 117
741 117
1 2 26 0 0 8320 0 37 29 0 0 3
607 110
607 105
741 105
1 3 25 0 0 0 0 50 28 0 0 2
765 117
896 117
1 1 26 0 0 0 0 29 28 0 0 2
765 105
896 105
0 0 27 0 0 8320 0 0 0 0 0 4
4 650
369 650
369 280
8 280
1 1 4 0 0 8320 0 32 30 0 0 4
317 642
317 705
405 705
405 715
2 1 4 0 0 0 0 32 31 0 0 3
326 642
326 695
405 695
2 1 28 0 0 4224 0 41 44 0 0 3
474 140
176 140
176 291
1 2 29 0 0 8320 0 43 40 0 0 3
166 291
166 120
474 120
2 1 5 0 0 8320 0 39 35 0 0 4
607 160
619 160
619 207
645 207
1 1 6 0 0 8320 0 39 36 0 0 4
607 150
632 150
632 190
645 190
1 1 30 0 0 8320 0 42 40 0 0 3
156 291
156 130
474 130
0 0 31 0 0 8320 0 0 0 0 0 6
470 90
470 80
610 80
610 200
470 200
470 90
82
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
630 60 726 104
634 64 722 96
22 4 CON.CABLE
P# 18777-
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
728 177 784 201
732 181 780 197
6 CONN.1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
768 150 784 174
772 154 780 170
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
769 137 785 161
773 141 781 157
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
768 124 784 148
772 128 780 144
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
768 114 784 138
772 118 780 134
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
768 101 784 125
772 105 780 121
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
767 89 783 113
771 93 779 109
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
819 90 851 114
823 94 847 110
3 RED
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
814 103 862 127
818 107 858 123
5 W/RED
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
821 139 869 163
825 143 865 159
5 W/GRN
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
821 152 853 176
825 156 849 172
3 GRN
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
167 311 191 375
171 315 187 363
9 D
I
R
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
147 311 171 375
151 315 167 363
9 +
5
V
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 17
158 311 182 415
162 315 178 395
17 P
U
L
S
E
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 26
142 501 222 565
146 505 218 553
26 CONVEYOR 
CONTROL
BOARD
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
120 297 152 321
124 301 148 317
3 TB2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
305 604 337 628
309 608 333 624
3 J11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
497 139 521 163
501 143 517 159
2 EN
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
497 129 529 153
501 133 525 149
3 DIR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
497 118 529 142
501 122 525 138
3 +5V
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
497 107 537 131
501 111 533 127
4 STEP
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
552 149 584 173
556 153 580 169
3 VDC
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
553 139 585 163
557 143 581 159
3 GND
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
560 128 584 152
564 132 580 148
2 A+
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
560 119 584 143
564 123 580 139
2 A-
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
560 109 584 133
564 113 580 129
2 B+
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
560 99 584 123
564 103 580 119
2 B-
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
494 77 590 101
498 81 586 97
11 STEP DRIVER
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
518 88 558 112
522 92 554 108
4 3535
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
324 346 356 370
328 350 352 366
3 TB4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
324 466 356 490
328 470 352 486
3 TB3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
227 606 259 630
231 610 255 626
3 PS1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
172 605 204 629
176 609 200 625
3 PS2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
118 605 150 629
122 609 146 625
3 PS3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
222 646 270 670
226 650 266 666
5 BOARD
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
222 659 278 683
226 663 274 679
6 AVAIL.
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
168 647 208 671
172 651 204 667
4 BUSY
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
115 647 155 671
119 651 151 667
4 SEND
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
9 647 57 671
13 651 53 667
5 PROX.
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
10 657 50 681
14 661 46 677
4 HIGH
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
58 647 106 671
62 651 102 667
5 PROX.
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
59 657 91 681
63 661 87 677
3 LOW
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
7 605 56 625
11 609 53 623
6 HI.LIM
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
56 605 105 625
60 609 102 623
6 LO.LIM
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 14
423 457 543 481
427 461 539 477
14 TERMINAL BLOCK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
750 414 766 438
754 418 762 434
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
750 404 766 428
754 408 762 424
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
675 426 707 450
679 430 703 446
3 YEL
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
676 415 708 439
680 419 704 435
3 PUR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
676 404 708 428
680 408 704 424
3 GRY
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
681 392 705 416
685 395 701 411
2 BL
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
944 440 960 464
948 444 956 460
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 15
889 452 1017 476
893 456 1013 472
15 (PCB UNLOADING)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
886 348 998 372
890 352 994 368
13 (PCB LOADING)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
944 337 960 361
948 341 956 357
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
673 289 697 313
677 292 693 308
2 BL
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
670 302 702 326
674 306 698 322
3 GRY
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
671 313 703 337
675 317 699 333
3 PUR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
670 325 702 349
674 329 698 345
3 YEL
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
746 289 762 313
750 293 758 309
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
747 300 763 324
751 304 759 320
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
747 314 763 338
751 318 759 334
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
750 391 766 415
754 395 762 411
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
747 325 763 349
751 329 759 345
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
750 429 766 453
754 433 762 449
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
747 339 763 363
751 343 759 359
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
747 351 763 375
751 355 759 371
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
749 442 765 466
753 446 761 462
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
749 455 765 479
753 459 761 475
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
791 288 815 312
795 292 811 308
2 LB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
786 301 818 325
790 305 814 321
3 GRY
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
786 313 818 337
790 317 814 333
3 BLK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
793 325 817 349
797 329 813 345
2 DB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
797 391 821 415
801 395 817 411
2 LB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
795 404 827 428
799 408 823 424
3 GRY
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
794 416 826 440
798 420 822 436
3 BLK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
797 428 821 452
801 432 817 448
2 DB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
710 478 766 502
714 482 762 498
6 CONN.3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
711 265 767 289
715 269 763 285
6 CONN.2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 30
681 529 929 553
685 533 925 549
30 * CONN.1,2&3 P#17028- & 17029-
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 23
480 283 672 307
484 287 668 303
23 4 CON.RIB.WIRE P#19210-
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
