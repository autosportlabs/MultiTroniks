CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
20 80 780 576
7 5.000 V
7 5.000 V
3 GND
1000 10
24 100 0 1 0
20 Package,Description,
61 C:\PROGRAM FILES\MICROCODE ENGINEERING\CIRCUITMAKER 6\BOM.DAT
0 7
20 80 780 576
143654930 0
0
0
0
0
0
0
34
7 Ground~
168 194 199 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8953 0 0
0
0
10 Capacitor~
219 194 175 0 2 5
0 2 9
0
0 0 576 90
15 .01uF CER. CAP.
-30 -5 75 3
2 C2
14 -15 28 -7
0
0
11 %D %1 %2 %V
0
0
7 CapCer1
5

0 1 2 1 2 -1610612704
67 0 0 0 1 0 0 0
1 C
4441 0 0
0
0
7 Ground~
168 487 177 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3618 0 0
0
0
7 Ground~
168 529 168 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6153 0 0
0
0
12 NPN Trans:C~
219 524 105 0 3 7
0 3 6 2
0
0 0 960 0
6 2N3904
22 -2 64 6
2 Q2
36 -12 50 -4
0
0
14 %D %1 %2 %3 %M
0
0
5 TO-39
7

0 1 2 3 1 2 3 -1610612700
81 0 0 0 1 0 0 0
1 Q
5394 0 0
0
0
7 Ground~
168 156 326 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7734 0 0
0
0
10 Capacitor~
219 177 262 0 2 5
0 2 13
0
0 0 576 0
14 18pf CER. CAP.
-50 -18 48 -10
2 C4
-8 -28 6 -20
0
0
11 %D %1 %2 %V
0
0
7 CapCer1
5

0 1 2 1 2 -1610612676
67 0 0 0 1 0 0 0
1 C
9914 0 0
0
0
10 Capacitor~
219 176 225 0 2 5
0 2 14
0
0 0 576 0
14 18pf CER. CAP.
-49 -18 49 -10
2 C3
-8 -28 6 -20
0
0
11 %D %1 %2 %V
0
0
7 CapCer1
5

0 1 2 1 2 -1610612676
67 0 0 0 1 0 0 0
1 C
3747 0 0
0
0
8 Crystal~
219 207 241 0 2 5
0 13 14
0
0 0 576 90
8 4.000MHZ
13 -5 69 3
3 XL1
-8 25 13 33
0
0
11 %D %1 %2 %S
0
32 alias:XCRYSTAL {FREQ=1E6 RS=540}
5 XTAL1
5

0 1 2 1 2 0
88 0 0 0 1 0 0 0
4 XTAL
3549 0 0
0
0
7 Ground~
168 86 329 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7931 0 0
0
0
7 Ground~
168 600 481 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9325 0 0
0
0
7 Ground~
168 394 446 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8903 0 0
0
0
4 LED~
171 446 282 0 2 2
10 17 16
0
0 0 624 0
15 RED LED 5MM/3MM
-76 -4 29 4
2 D1
-24 4 -10 12
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3834 0 0
0
0
7 Ground~
168 446 444 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3363 0 0
0
0
12 NPN Trans:C~
219 441 370 0 3 7
0 16 5 2
0
0 0 832 0
6 2N3904
14 9 56 17
2 Q1
28 -1 42 7
0
0
14 %D %1 %2 %3 %M
0
0
5 TO-39
7

0 1 2 3 1 2 3 -1610612704
81 0 0 0 1 1 0 0
1 Q
7668 0 0
0
0
7 Ground~
168 93 208 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4718 0 0
0
0
7 Ground~
168 564 250 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3874 0 0
0
0
10 Polar Cap~
219 94 176 0 2 5
0 9 2
0
0 0 576 270
15 10uF ELEC. CAPA
-31 -1 74 7
2 C1
14 -11 28 -3
0
0
11 %D %1 %2 %V
0
0
7 CapPol1
5

0 1 2 1 2 -1610612720
67 0 0 0 1 0 0 0
1 C
6671 0 0
0
0
7 Ground~
168 381 219 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3789 0 0
0
0
4 CON2
94 59 61 0 2 5
0 11 3
4 CON2
1 0 4608 0
15 HEADER 2 PIN MO
-56 -30 49 -22
2 J1
-11 -40 3 -32
0
0
0
0
0
6 MOLEX2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 J
4871 0 0
0
0
4 CON2
94 594 61 0 2 5
0 11 3
4 CON2
2 0 4608 512
15 HEADER 2 PIN MO
-56 -30 49 -22
2 J2
-11 -40 3 -32
0
0
0
0
0
6 MOLEX2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 J
3750 0 0
0
0
4 CON3
94 679 429 0 3 7
0 2 16 7
4 CON3
3 0 4608 0
15 HEADER 3 PIN MO
-48 -31 57 -23
2 J3
-3 -41 11 -33
0
0
0
0
0
6 MOLEX3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 J
8778 0 0
0
0
4 CON3
94 677 295 0 3 7
0 10 8 15
4 CON3
4 0 4608 0
2 TP
-3 -31 11 -23
3 TP1
-6 -41 15 -33
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 J
538 0 0
0
0
8 PIC12671
94 334 254 0 8 17
0 14 13 4 15 10 8 2 9
8 PIC12671
5 0 6784 0
8 PIC12671
-49 -76 7 -68
2 U1
-28 -86 -14 -78
0
0
0
0
0
4 DIP8
17

0 2 3 4 5 6 7 8 1 2
3 4 5 6 7 8 1 -1610612720
0 0 0 0 1 1 0 0
1 U
6843 0 0
0
0
3 REG
94 566 191 0 3 7
0 12 2 9
3 REG
6 0 6912 512
13 5V REG  78L05
-46 -14 45 -6
2 Q3
-5 -24 9 -16
0
0
0
0
0
5 TO-39
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 Q
3136 0 0
0
0
6 VACSEN
94 63 269 0 6 13
0 95 9 8 2 96 97
6 VACSEN
7 0 2560 90
15 PRESSURE SENSOR
-54 -30 51 -22
2 S1
-8 -40 6 -32
0
0
0
0
0
7 VAC SEN
13

0 1 2 3 4 5 6 1 2 3
4 5 6 0
0 0 0 512 1 0 0 0
1 J
5950 0 0
0
0
9 Resistor~
219 487 138 0 4 5
0 6 2 0 -1
0
0 0 864 270
3 47k
7 0 28 8
2 R7
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612676
82 0 0 0 1 0 0 0
1 R
5670 0 0
0
0
9 Resistor~
219 462 105 0 2 5
0 10 6
0
0 0 864 0
4 2.2k
-14 -14 14 -6
2 R6
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612671
82 0 0 0 1 0 0 0
1 R
6828 0 0
0
0
9 Resistor~
219 145 102 0 2 5
0 4 3
0
0 0 864 90
4 750k
8 0 36 8
2 R5
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612720
82 0 0 0 1 0 0 0
1 R
6735 0 0
0
0
9 Resistor~
219 227 243 0 2 5
0 13 14
0
0 0 864 90
3 10M
5 0 26 8
2 R1
7 -10 21 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612676
82 0 0 0 1 0 0 0
1 R
8365 0 0
0
0
9 Resistor~
219 446 238 0 2 5
0 17 9
0
0 0 864 90
3 470
5 -5 26 3
2 R4
8 -15 22 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612720
82 0 0 0 1 0 0 0
1 R
4132 0 0
0
0
9 Resistor~
219 394 336 0 2 5
0 5 15
0
0 0 864 90
3 10k
5 -5 26 3
2 R2
8 -15 22 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612720
82 0 0 0 1 0 0 0
1 R
4551 0 0
0
0
9 Resistor~
219 394 405 0 4 5
0 5 2 0 -1
0
0 0 864 270
3 47k
7 0 28 8
2 R3
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612676
82 0 0 0 1 0 0 0
1 R
3635 0 0
0
0
9 Resistor~
219 628 351 0 2 5
0 7 12
0
0 0 864 90
7 1K/0.5W
1 -4 50 4
2 R8
8 -15 22 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612676
82 0 0 0 1 0 0 0
1 R
3973 0 0
0
0
43
1 0 3 0 0 4096 0 5 0 0 19 2
529 87
529 61
2 0 3 0 0 0 0 29 0 0 19 2
145 84
145 61
1 3 4 0 0 4224 0 29 24 0 0 3
145 120
145 288
257 288
2 1 2 0 0 4096 0 33 12 0 0 2
394 423
394 440
0 1 5 0 0 4096 0 0 32 35 0 2
394 370
394 354
2 1 2 0 0 0 0 27 3 0 0 2
487 156
487 171
1 0 6 0 0 4096 0 27 0 0 17 2
487 120
487 105
1 3 7 0 0 4224 0 34 22 0 0 3
628 369
628 438
673 438
1 1 2 0 0 4224 0 22 11 0 0 3
673 418
600 418
600 475
3 0 8 0 0 12416 0 26 0 0 11 4
70 289
112 289
112 472
381 472
6 2 8 0 0 0 0 24 23 0 0 6
369 244
381 244
381 472
498 472
498 294
671 294
1 1 2 0 0 0 0 2 1 0 0 2
194 184
194 193
2 0 9 0 0 4096 0 2 0 0 43 2
194 166
194 143
0 1 10 0 0 4096 0 0 23 16 0 4
429 266
589 266
589 284
671 284
2 1 2 0 0 0 0 25 17 0 0 2
564 225
564 244
1 5 10 0 0 8320 0 28 24 0 0 4
444 105
429 105
429 274
369 274
2 2 6 0 0 4224 0 28 5 0 0 2
480 105
506 105
3 1 2 0 0 0 0 5 4 0 0 2
529 123
529 162
2 2 3 0 0 4224 0 20 21 0 0 2
66 61
573 61
1 1 11 0 0 4224 0 20 21 0 0 2
66 51
573 51
3 0 9 0 0 4096 0 25 0 0 40 2
527 203
446 203
1 2 12 0 0 8320 0 25 34 0 0 3
601 202
628 202
628 333
1 0 13 0 0 4096 0 9 0 0 29 2
207 252
207 262
2 0 14 0 0 4096 0 9 0 0 30 2
207 230
207 225
1 2 13 0 0 8192 0 30 24 0 0 5
227 261
227 262
242 262
242 258
257 258
1 2 14 0 0 4096 0 24 30 0 0 4
256 227
240 227
240 225
227 225
0 1 2 0 0 0 0 0 6 28 0 2
156 262
156 320
1 1 2 0 0 0 0 8 7 0 0 4
167 225
156 225
156 262
168 262
2 1 13 0 0 4224 0 7 30 0 0 3
186 262
227 262
227 261
2 2 14 0 0 4224 0 8 30 0 0 2
185 225
227 225
4 1 2 0 0 0 0 26 10 0 0 3
70 279
86 279
86 323
2 0 9 0 0 8192 0 26 0 0 43 3
70 299
126 299
126 143
0 3 15 0 0 4224 0 0 23 36 0 2
393 304
671 304
0 2 16 0 0 4224 0 0 22 38 0 4
446 325
569 325
569 428
673 428
2 1 5 0 0 4224 0 15 33 0 0 3
423 370
394 370
394 387
4 2 15 0 0 0 0 24 32 0 0 3
370 304
394 304
394 318
3 1 2 0 0 0 0 15 14 0 0 2
446 388
446 438
2 1 16 0 0 0 0 13 15 0 0 2
446 292
446 352
1 1 17 0 0 4224 0 31 13 0 0 2
446 256
446 272
0 2 9 0 0 4224 0 0 31 43 0 3
253 143
446 143
446 220
7 1 2 0 0 0 0 24 19 0 0 3
371 204
381 204
381 213
2 1 2 0 0 0 0 18 16 0 0 2
93 183
93 202
1 8 9 0 0 0 0 18 24 0 0 5
93 166
93 143
253 143
253 204
258 204
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
