CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 800 30 80 9
0 66 800 569
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
61 C:\PROGRAM FILES\MICROCODE ENGINEERING\CIRCUITMAKER 6\BOM.DAT
0 7
0 66 800 569
146341906 0
0
6 Title:
5 Name:
10 09-17-1998
0
0
85
11 SPDT Relay~
176 894 694 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 4192 512
7 12VSPDT
-25 -35 24 -27
4 RLY3
-14 -45 14 -37
0
0
20 %D %1 %2 %3 %4 %5 %S
0
45 alias:XSPDTRELAY {PULLIN=9.6 RESISTANCE=1000}
4 DIP4
11

0 1 2 3 4 5 1 2 3 4
5 0
88 0 0 0 0 0 0 0
3 RLY
8953 0 0
0
0
10 Capacitor~
219 609 1147 0 2 5
0 2 3
0
0 0 832 90
3 1uF
11 0 32 8
3 C12
11 -10 32 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -1610612676
67 0 0 0 1 0 0 0
1 C
4441 0 0
0
0
7 Ground~
168 457 1205 0 1 3
0 2
0
0 0 53344 0
0
5 GND14
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3618 0 0
0
0
7 Ground~
168 285 1241 0 1 3
0 2
0
0 0 53344 0
0
5 GND13
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6153 0 0
0
0
10 Capacitor~
219 236 1165 0 2 5
0 2 13
0
0 0 832 90
3 1uF
11 0 32 8
3 C11
11 -10 32 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -1610612676
67 0 0 0 1 0 0 0
1 C
5394 0 0
0
0
7 Ground~
168 604 1086 0 1 3
0 2
0
0 0 53344 0
0
5 GND12
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7734 0 0
0
0
10 Capacitor~
219 784 913 0 2 5
0 2 3
0
0 0 832 90
3 1uF
11 0 32 8
3 C10
11 -10 32 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -1610612720
67 0 0 0 1 0 0 0
1 C
9914 0 0
0
0
10 Capacitor~
219 619 950 0 2 5
0 2 3
0
0 0 832 90
3 1uF
8 1 29 9
2 C9
9 -14 23 -6
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -1610612720
67 0 0 0 1 0 0 0
1 C
3747 0 0
0
0
6 Diode~
219 946 712 0 2 5
0 37 15
0
0 0 64 0
5 DIODE
-18 -18 17 -10
3 D43
-11 -28 10 -20
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
3549 0 0
0
0
6 Diode~
219 757 727 0 2 5
0 33 15
0
0 0 64 0
5 DIODE
-18 -18 17 -10
3 D42
-11 -28 10 -20
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
7931 0 0
0
0
6 Diode~
219 590 753 0 2 5
0 36 15
0
0 0 64 0
5 DIODE
-18 -18 17 -10
3 D41
-11 -28 10 -20
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
9325 0 0
0
0
7 Ground~
168 848 694 0 1 3
0 2
0
0 0 53344 0
0
5 GND11
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8903 0 0
0
0
7 Ground~
168 652 713 0 1 3
0 2
0
0 0 53344 0
0
5 GND10
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3834 0 0
0
0
7 Ground~
168 473 741 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3363 0 0
0
0
11 Contacts:A~
214 893 654 0 10 11
0 2 34 35 0 0 0 0 0 0
1
0
0 0 96 512
6 NORMAL
-23 -17 19 -9
4 RLY5
-16 -27 12 -19
0
0
17 %D %1 %2 %3 %I %S
0
15 alias:XCONTACTS
4 SIP3
7

0 1 2 3 1 2 3 0
88 0 0 0 1 0 0 0
3 RLY
7668 0 0
0
0
11 Contacts:A~
214 893 630 0 10 11
0 30 164 33 0 0 0 0 0 0
1
0
0 0 96 512
6 NORMAL
-23 -17 19 -9
4 RLY6
-16 -27 12 -19
0
0
17 %D %1 %2 %3 %I %S
0
15 alias:XCONTACTS
4 SIP3
7

0 1 2 3 1 2 3 0
88 0 0 512 1 0 0 0
3 RLY
4718 0 0
0
0
11 SPDT Relay~
176 700 708 0 10 11
0 2 165 31 15 33 0 0 0 0
1
0
0 0 4192 512
7 12VSPDT
-27 -35 22 -27
4 RLY2
-16 -45 12 -37
0
0
20 %D %1 %2 %3 %4 %5 %S
0
45 alias:XSPDTRELAY {PULLIN=9.6 RESISTANCE=1000}
4 DIP4
11

0 1 2 3 4 5 1 2 3 4
5 0
88 0 0 512 1 0 0 0
3 RLY
3874 0 0
0
0
11 Contacts:A~
214 698 668 0 10 11
0 2 6 32 0 0 0 0 0 0
1
0
0 0 96 512
6 NORMAL
-23 -17 19 -9
4 RLY4
-16 -27 12 -19
0
0
17 %D %1 %2 %3 %I %S
0
15 alias:XCONTACTS
4 SIP3
7

0 1 2 3 1 2 3 0
88 0 0 0 1 0 0 0
3 RLY
6671 0 0
0
0
11 SPDT Relay~
176 534 733 0 10 11
0 2 38 36 15 36 0 0 0 0
1
0
0 0 2144 512
7 12VSPDT
-27 -35 22 -27
4 RLY1
-16 -45 12 -37
0
0
20 %D %1 %2 %3 %4 %5 %S
0
45 alias:XSPDTRELAY {PULLIN=9.6 RESISTANCE=1000}
4 DIP4
11

0 1 2 3 4 5 1 2 3 4
5 0
88 0 0 0 1 1 0 0
3 RLY
3789 0 0
0
0
6 74-244
94 691 253 0 20 41
0 154 153 152 151 150 149 148 147 2
2 2 106 107 108 109 111 112 113 114
22
6 74-244
1 0 15232 0
5 74244
-18 -64 17 -56
2 U3
-7 -74 7 -66
0
0
0
0
0
5 DIP20
41

0 2 17 4 15 6 13 8 11 1
19 10 9 12 7 14 5 16 3 18
20 2 17 4 15 6 13 8 11 1
19 10 9 12 7 14 5 16 3 18
20 0
0 0 0 0 1 0 0 0
1 U
4871 0 0
0
0
6 26LS32
94 412 590 0 16 33
0 46 45 40 166 39 44 43 2 50
49 42 2 41 48 47 3
6 26LS32
2 0 6816 0
0
2 U7
-7 -55 7 -47
0
0
0
0
0
5 DIP16
33

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 1 2 3
4 5 6 7 8 9 10 11 12 13
14 15 16 0
0 0 0 512 1 0 0 0
1 U
3750 0 0
0
0
6 74-244
94 692 524 0 20 41
0 138 137 136 135 134 133 132 131 2
2 2 74 75 76 77 79 80 81 82
22
6 74-244
4 0 15232 0
5 74244
-18 -64 17 -56
2 U5
-7 -74 7 -66
0
0
0
0
0
5 DIP20
41

0 2 17 4 15 6 13 8 11 1
19 10 9 12 7 14 5 16 3 18
20 2 17 4 15 6 13 8 11 1
19 10 9 12 7 14 5 16 3 18
20 0
0 0 0 0 1 0 0 0
1 U
8778 0 0
0
0
6 74-244
94 584 403 0 20 41
0 146 145 144 143 142 141 140 139 2
2 2 90 91 92 93 95 96 97 98
22
6 74-244
5 0 15232 0
5 74244
-18 -64 17 -56
2 U4
-7 -74 7 -66
0
0
0
0
0
5 DIP20
41

0 2 17 4 15 6 13 8 11 1
19 10 9 12 7 14 5 16 3 18
20 2 17 4 15 6 13 8 11 1
19 10 9 12 7 14 5 16 3 18
20 0
0 0 0 0 1 0 0 0
1 U
538 0 0
0
0
6 74-244
94 579 123 0 20 41
0 162 161 160 159 158 157 156 155 2
2 2 122 123 124 125 127 128 129 130
22
6 74-244
6 0 15232 0
5 74244
-18 -64 17 -56
2 U2
-7 -74 7 -66
0
0
0
0
0
5 DIP20
41

0 2 17 4 15 6 13 8 11 1
19 10 9 12 7 14 5 16 3 18
20 2 17 4 15 6 13 8 11 1
19 10 9 12 7 14 5 16 3 18
20 0
0 0 0 0 1 0 0 0
1 U
6843 0 0
0
0
6 CON-64
94 339 305 0 129 129
0 15 2 22 20 21 23 25 26 11
27 28 16 17 18 19 31 32 34 35
38 43 44 39 40 45 46 47 48 41
42 49 50 131 132 133 134 135 136 137
138 139 140 141 142 143 144 145 146 147
148 149 150 151 152 153 154 155 156 157
158 159 160 161 162 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 -1610612212
6 CON-64
7 0 4736 0
0
2 J2
0 -163 14 -155
0
0
0
0
0
0
129

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 21 22 23 24 25 26 27 28 29
30 31 32 33 34 35 36 37 38 39
40 41 42 43 44 45 46 47 48 49
50 51 52 53 54 55 56 57 58 59
60 61 62 63 64 1 2 3 4 5
6 7 8 9 10 11 12 13 14 15
16 17 18 19 20 21 22 23 24 25
26 27 28 29 30 31 32 33 34 35
36 37 38 39 40 41 42 43 44 45
46 47 48 49 50 51 52 53 54 55
56 57 58 59 60 61 62 63 64 0
0 0 0 0 1 0 0 0
1 J
3136 0 0
0
0
7 Ground~
168 648 598 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5950 0 0
0
0
7 Ground~
168 533 475 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5670 0 0
0
0
7 Ground~
168 650 328 0 1 3
0 2
0
0 0 53344 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6828 0 0
0
0
7 Ground~
168 533 200 0 1 3
0 2
0
0 0 53344 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6735 0 0
0
0
4 LED~
171 890 70 0 2 2
10 130 126
0
0 0 112 90
4 LED1
-12 -21 16 -13
2 D1
-5 -31 9 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
8365 0 0
0
0
4 LED~
171 870 86 0 2 2
10 129 121
0
0 0 112 90
4 LED1
-12 -21 16 -13
2 D2
-5 -31 9 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
4132 0 0
0
0
4 LED~
171 890 102 0 2 2
10 128 120
0
0 0 112 90
4 LED1
-12 -21 16 -13
2 D3
-5 -31 9 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
4551 0 0
0
0
4 LED~
171 869 117 0 2 2
10 127 119
0
0 0 112 90
4 LED1
-12 -21 16 -13
2 D4
-5 -31 9 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3635 0 0
0
0
7 RSIP10~
219 1021 110 0 10 21
0 2 168 126 121 120 119 118 117 116
115
0
0 0 832 270
2 1k
-9 -52 5 -44
2 R1
-9 -62 5 -54
0
0
125 %DA %1 %2 %V
%DB %1 %3 %V
%DC %1 %4 %V
%DD %1 %5 %V
%DE %1 %6 %V
%DF %1 %7 %V
%DG %1 %8 %V
%DH %1 %9 %V
%DI %1 %10 %V
0
0
5 SIP10
21

0 1 2 3 4 5 6 7 8 9
10 1 2 3 4 5 6 7 8 9
10 0
82 0 0 512 1 0 0 0
1 R
3973 0 0
0
0
4 LED~
171 866 178 0 2 2
10 122 115
0
0 0 112 90
4 LED1
-12 -21 16 -13
2 D5
-5 -31 9 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3851 0 0
0
0
4 LED~
171 886 163 0 2 2
10 123 116
0
0 0 112 90
4 LED1
-12 -21 16 -13
2 D6
-5 -31 9 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
8383 0 0
0
0
4 LED~
171 869 148 0 2 2
10 124 117
0
0 0 112 90
4 LED1
-12 -21 16 -13
2 D7
-5 -31 9 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
9334 0 0
0
0
4 LED~
171 889 131 0 2 2
10 125 118
0
0 0 112 90
4 LED1
-12 -21 16 -13
2 D8
-5 -31 9 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
7471 0 0
0
0
4 LED~
171 886 260 0 2 2
10 109 102
0
0 0 112 90
4 LED1
-12 -21 16 -13
2 D9
-5 -31 9 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3334 0 0
0
0
4 LED~
171 866 276 0 2 2
10 108 101
0
0 0 112 90
4 LED1
-12 -21 16 -13
3 D10
-8 -31 13 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3559 0 0
0
0
4 LED~
171 886 292 0 2 2
10 107 100
0
0 0 112 90
4 LED1
-12 -21 16 -13
3 D11
-8 -31 13 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
984 0 0
0
0
4 LED~
171 866 307 0 2 2
10 106 99
0
0 0 112 90
4 LED1
-12 -21 16 -13
3 D12
-8 -31 13 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
7557 0 0
0
0
7 RSIP10~
219 1021 264 0 10 21
0 2 169 110 105 104 103 102 101 100
99
0
0 0 832 270
2 1k
-9 -52 5 -44
2 R2
-9 -62 5 -54
0
0
125 %DA %1 %2 %V
%DB %1 %3 %V
%DC %1 %4 %V
%DD %1 %5 %V
%DE %1 %6 %V
%DF %1 %7 %V
%DG %1 %8 %V
%DH %1 %9 %V
%DI %1 %10 %V
0
0
5 SIP10
21

0 1 2 3 4 5 6 7 8 9
10 1 2 3 4 5 6 7 8 9
10 0
82 0 0 512 1 0 0 0
1 R
3146 0 0
0
0
4 LED~
171 868 243 0 2 2
10 111 103
0
0 0 112 90
4 LED1
-12 -21 16 -13
3 D13
-8 -31 13 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
5687 0 0
0
0
4 LED~
171 885 227 0 2 2
10 112 104
0
0 0 112 90
4 LED1
-12 -21 16 -13
3 D14
-8 -31 13 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
7939 0 0
0
0
4 LED~
171 867 211 0 2 2
10 113 105
0
0 0 112 90
4 LED1
-12 -21 16 -13
3 D15
-8 -31 13 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3308 0 0
0
0
4 LED~
171 885 195 0 2 2
10 114 110
0
0 0 112 90
4 LED1
-12 -21 16 -13
3 D16
-8 -31 13 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3408 0 0
0
0
4 LED~
171 885 393 0 2 2
10 93 86
0
0 0 112 90
4 LED1
-12 -21 16 -13
3 D17
-8 -31 13 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
9773 0 0
0
0
4 LED~
171 866 407 0 2 2
10 92 85
0
0 0 112 90
4 LED1
-12 -21 16 -13
3 D18
-8 -31 13 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
691 0 0
0
0
4 LED~
171 885 422 0 2 2
10 91 84
0
0 0 112 90
4 LED1
-12 -21 16 -13
3 D19
-8 -31 13 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
7834 0 0
0
0
4 LED~
171 865 438 0 2 2
10 90 83
0
0 0 112 90
4 LED1
-12 -21 16 -13
3 D20
-8 -31 13 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3588 0 0
0
0
7 RSIP10~
219 1019 395 0 10 21
0 2 170 94 89 88 87 86 85 84
83
0
0 0 832 270
2 1k
-9 -52 5 -44
2 R3
-9 -62 5 -54
0
0
125 %DA %1 %2 %V
%DB %1 %3 %V
%DC %1 %4 %V
%DD %1 %5 %V
%DE %1 %6 %V
%DF %1 %7 %V
%DG %1 %8 %V
%DH %1 %9 %V
%DI %1 %10 %V
0
0
5 SIP10
21

0 1 2 3 4 5 6 7 8 9
10 1 2 3 4 5 6 7 8 9
10 0
82 0 0 512 1 0 0 0
1 R
4528 0 0
0
0
4 LED~
171 866 378 0 2 2
10 95 87
0
0 0 112 90
4 LED1
-12 -21 16 -13
3 D21
-8 -31 13 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3303 0 0
0
0
4 LED~
171 885 363 0 2 2
10 96 88
0
0 0 112 90
4 LED1
-12 -21 16 -13
3 D22
-8 -31 13 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
9654 0 0
0
0
4 LED~
171 867 347 0 2 2
10 97 89
0
0 0 112 90
4 LED1
-12 -21 16 -13
3 D23
-8 -31 13 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
9791 0 0
0
0
4 LED~
171 885 330 0 2 2
10 98 94
0
0 0 112 90
4 LED1
-12 -21 16 -13
3 D24
-8 -31 13 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
4589 0 0
0
0
4 LED~
171 864 523 0 2 2
10 77 70
0
0 0 112 90
4 LED1
-12 -21 16 -13
3 D25
-8 -31 13 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
964 0 0
0
0
4 LED~
171 888 541 0 2 2
10 76 69
0
0 0 112 90
4 LED1
-12 -21 16 -13
3 D26
-8 -31 13 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
9151 0 0
0
0
4 LED~
171 865 555 0 2 2
10 75 68
0
0 0 112 90
4 LED1
-12 -21 16 -13
3 D27
-8 -31 13 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
4745 0 0
0
0
4 LED~
171 887 571 0 2 2
10 74 67
0
0 0 112 90
4 LED1
-12 -21 16 -13
3 D28
-8 -31 13 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
8433 0 0
0
0
7 RSIP10~
219 1019 528 0 10 21
0 2 171 78 73 72 71 70 69 68
67
0
0 0 832 270
2 1k
-9 -52 5 -44
2 R4
-9 -62 5 -54
0
0
125 %DA %1 %2 %V
%DB %1 %3 %V
%DC %1 %4 %V
%DD %1 %5 %V
%DE %1 %6 %V
%DF %1 %7 %V
%DG %1 %8 %V
%DH %1 %9 %V
%DI %1 %10 %V
0
0
5 SIP10
21

0 1 2 3 4 5 6 7 8 9
10 1 2 3 4 5 6 7 8 9
10 0
82 0 0 512 1 0 0 0
1 R
4221 0 0
0
0
4 LED~
171 887 510 0 2 2
10 79 71
0
0 0 112 90
4 LED1
-12 -21 16 -13
3 D29
-8 -31 13 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
8348 0 0
0
0
4 LED~
171 864 496 0 2 2
10 80 72
0
0 0 112 90
4 LED1
-12 -21 16 -13
3 D30
-8 -31 13 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
5299 0 0
0
0
4 LED~
171 886 481 0 2 2
10 81 73
0
0 0 112 90
4 LED1
-12 -21 16 -13
3 D31
-8 -31 13 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
7393 0 0
0
0
4 LED~
171 864 465 0 2 2
10 82 78
0
0 0 112 90
4 LED1
-12 -21 16 -13
3 D32
-8 -31 13 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
6917 0 0
0
0
7 Ground~
168 985 587 0 1 3
0 2
0
0 0 53344 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8767 0 0
0
0
7 Ground~
168 238 153 0 1 3
0 2
0
0 0 53344 0
0
4 GND8
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3606 0 0
0
0
10 Polar Cap~
219 239 115 0 2 5
0 22 2
0
0 0 832 270
9 220uF/16V
-73 1 -10 9
2 C1
-26 -10 -12 -2
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
6970 0 0
0
0
10 Capacitor~
219 279 113 0 2 5
0 2 22
0
0 0 832 90
5 0.1uF
21 1 56 9
2 C2
23 -10 37 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
343 0 0
0
0
10 Capacitor~
219 651 173 0 2 5
0 2 22
0
0 0 832 90
3 1uF
11 0 32 8
2 C3
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7197 0 0
0
0
10 Capacitor~
219 763 306 0 2 5
0 2 22
0
0 0 832 90
3 1uF
11 0 32 8
2 C4
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3623 0 0
0
0
10 Capacitor~
219 649 456 0 2 5
0 2 22
0
0 0 832 90
3 1uF
11 0 32 8
2 C5
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7656 0 0
0
0
10 Capacitor~
219 753 575 0 2 5
0 2 22
0
0 0 832 90
3 1uF
11 0 32 8
2 C6
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
5365 0 0
0
0
7 Ground~
168 307 663 0 1 3
0 2
0
0 0 53344 0
0
4 GND9
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4557 0 0
0
0
10 Capacitor~
219 532 587 0 2 5
0 2 3
0
0 0 832 90
3 1uF
11 0 32 8
2 C8
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3489 0 0
0
0
4 2003
94 934 889 0 16 33
0 4 173 8 20 174 175 12 2 30
176 7 21 11 27 28 15
4 2003
8 0 6784 0
0
2 U1
-7 -56 7 -48
0
0
0
0
0
0
33

0 1 2 3 4 5 6 7 8 16
15 14 13 12 11 10 9 1 2 3
4 5 6 7 8 16 15 14 13 12
11 10 9 0
0 0 0 512 1 1 0 0
1 U
345 0 0
0
0
6 74-138
94 573 895 0 16 33
0 19 18 17 16 16 3 177 2 178
29 179 180 181 182 183 3
6 74-138
9 0 4864 0
5 74138
-18 -42 17 -34
2 U8
-7 -55 7 -47
0
0
0
0
0
5 DIP16
33

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 1 2 3
4 5 6 7 8 9 10 11 12 13
14 15 16 -1610612708
0 0 0 512 1 0 0 0
1 U
3374 0 0
0
0
5 74-00
94 720 899 0 14 29
0 29 29 4 26 25 24 2 23 24
24 184 185 186 3
5 74-00
10 0 4864 0
4 7400
-15 -31 13 -23
2 U9
-7 -47 7 -39
0
0
0
0
0
0
29

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 1 2 3 4 5
6 7 8 9 10 11 12 13 14 0
0 0 0 512 1 0 0 0
1 U
5866 0 0
0
0
5 74-00
94 531 1128 0 14 29
0 10 10 8 6 6 5 2 216 217
218 9 8 8 3
5 74-00
12 0 4736 0
0
3 U10
-11 -47 10 -39
0
0
0
0
0
0
29

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 1 2 3 4 5
6 7 8 9 10 11 12 13 14 0
0 0 0 512 1 0 0 0
0
631 0 0
0
0
9 Resistor~
219 883 951 0 2 5
0 11 12
0
0 0 864 90
2 1k
11 0 25 8
3 R11
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612604
82 0 0 0 1 0 0 0
1 R
745 0 0
0
0
9 Resistor~
219 334 1174 0 3 5
0 2 10 -1
0
0 0 864 90
2 1k
11 0 25 8
3 R10
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612700
82 0 0 0 1 0 0 0
1 R
7222 0 0
0
0
9 Resistor~
219 286 1115 0 2 5
0 13 10
0
0 0 864 0
2 1k
-7 -14 7 -6
2 R9
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612704
82 0 0 0 1 0 0 0
1 R
4508 0 0
0
0
9 Resistor~
219 236 1054 0 2 5
0 14 13
0
0 0 864 270
2 1k
8 0 22 8
2 R8
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612676
82 0 0 0 1 0 0 0
1 R
3738 0 0
0
0
9 Resistor~
219 864 951 0 3 5
0 2 12 -1
0
0 0 864 90
2 1k
8 0 22 8
2 R7
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612604
82 0 0 0 1 0 0 0
1 R
91 0 0
0
0
9 Resistor~
219 724 622 0 2 5
0 34 3
0
0 0 864 180
2 1k
6 8 20 16
2 R6
-16 8 -2 16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612720
82 0 0 0 1 0 0 0
1 R
4965 0 0
0
0
225
30 0 0 0 0 0 0 25 0 0 5 3
313 431
299 431
299 440
1 0 0 0 0 0 0 25 0 0 57 2
313 170
279 170
0 0 0 0 0 0 0 0 0 109 4 3
307 626
306 626
306 485
32 33 0 0 0 0 0 25 25 0 0 6
313 449
306 449
306 485
385 485
385 449
379 449
0 31 0 0 0 0 0 0 25 6 0 7
997 921
997 1025
440 1025
440 911
268 911
268 440
313 440
0 16 0 0 0 0 0 0 76 92 0 3
997 752
997 923
965 923
11 29 0 0 0 0 0 76 25 0 0 8
965 873
1044 873
1044 1239
373 1239
373 985
256 985
256 422
313 422
28 11 0 0 0 0 0 25 79 0 0 8
313 413
246 413
246 975
383 975
383 1229
591 1229
591 1137
564 1137
27 1 0 0 0 0 0 25 83 0 0 3
313 404
236 404
236 1036
2 0 0 0 0 0 0 5 0 0 47 2
236 1156
236 1115
0 0 0 0 0 0 0 0 0 12 21 2
488 1115
335 1115
2 1 0 0 0 0 0 79 79 0 0 4
498 1119
488 1119
488 1110
498 1110
10 0 0 0 0 0 0 77 0 0 78 4
606 922
639 922
639 886
675 886
2 0 0 0 0 0 0 8 0 0 77 2
619 941
619 867
0 3 0 0 0 0 0 0 16 16 0 3
730 727
730 637
879 637
1 5 0 0 0 0 0 10 17 0 0 2
747 727
714 727
0 2 0 0 0 0 0 0 85 108 0 6
533 563
619 563
619 623
619 623
619 622
706 622
1 0 0 0 0 0 0 1 0 0 96 2
878 676
847 676
0 7 0 0 0 0 0 0 22 79 0 5
793 852
793 612
633 612
633 542
659 542
6 6 0 0 0 0 0 79 22 0 0 4
498 1155
345 1155
345 533
659 533
0 5 0 0 0 0 0 0 22 46 0 3
335 1115
335 524
659 524
4 0 0 0 0 0 0 22 0 0 102 2
659 515
199 515
3 0 0 0 0 0 0 22 0 0 104 2
659 506
209 506
2 0 0 0 0 0 0 22 0 0 28 2
659 497
492 497
1 0 0 0 0 0 0 22 0 0 29 2
659 488
502 488
15 35 0 0 0 0 0 21 25 0 0 6
445 572
473 572
473 487
409 487
409 431
379 431
14 36 0 0 0 0 0 21 25 0 0 6
445 581
482 581
482 477
419 477
419 422
379 422
13 37 0 0 0 0 0 21 25 0 0 6
445 590
492 590
492 467
429 467
429 413
379 413
11 38 0 0 0 0 0 21 25 0 0 6
445 608
502 608
502 457
438 457
438 404
379 404
10 39 0 0 0 0 0 21 25 0 0 6
445 617
511 617
511 448
449 448
449 395
379 395
9 40 0 0 0 0 0 21 25 0 0 6
445 626
520 626
520 439
459 439
459 386
379 386
1 0 2 0 0 8192 0 2 0 0 34 3
609 1156
609 1191
458 1191
2 0 3 0 0 4096 0 2 0 0 35 2
609 1138
609 1110
7 1 2 0 0 0 0 79 3 0 0 4
498 1164
458 1164
458 1199
457 1199
0 14 3 0 0 12288 0 0 79 77 0 4
783 839
837 839
837 1110
564 1110
0 0 3 0 0 0 0 0 0 77 17 2
619 839
619 623
0 2 6 0 0 12416 0 0 18 38 0 5
487 1146
487 1145
361 1145
361 661
684 661
5 4 6 0 0 0 0 79 79 0 0 4
498 1146
487 1146
487 1137
498 1137
0 3 8 0 0 4224 0 0 76 41 0 4
588 1102
848 1102
848 873
902 873
0 12 8 0 0 0 0 0 79 41 0 3
575 1123
575 1128
564 1128
3 13 8 0 0 0 0 79 79 0 0 8
498 1128
467 1128
467 1080
588 1080
588 1123
575 1123
575 1119
564 1119
1 0 11 0 0 4096 0 80 0 0 64 2
883 969
883 1053
2 0 12 0 0 4096 0 80 0 0 68 2
883 933
883 913
1 0 2 0 0 0 0 4 0 0 45 2
285 1235
285 1205
1 1 2 0 0 0 0 5 81 0 0 4
236 1174
236 1205
334 1205
334 1192
2 2 10 0 0 0 0 82 81 0 0 5
304 1115
335 1115
335 1115
334 1115
334 1156
2 1 13 0 0 4224 0 83 82 0 0 3
236 1072
236 1115
268 1115
0 2 2 0 0 0 0 0 68 57 0 2
238 138
238 122
0 1 2 0 0 0 0 0 69 57 0 2
279 139
279 122
0 12 16 0 0 16512 0 0 25 70 0 6
532 899
476 899
476 868
97 868
97 269
313 269
3 13 17 0 0 16512 0 77 25 0 0 6
540 886
485 886
485 856
106 856
106 278
313 278
2 14 18 0 0 16512 0 77 25 0 0 6
540 877
494 877
494 846
115 846
115 287
313 287
1 15 19 0 0 16512 0 77 25 0 0 7
540 868
503 868
503 835
124 835
124 297
313 297
313 296
4 4 20 0 0 24704 0 76 25 0 0 8
902 883
909 883
909 1071
391 1071
391 964
12 964
12 197
313 197
5 12 21 0 0 8320 0 25 76 0 0 8
313 206
23 206
23 952
400 952
400 1062
1035 1062
1035 883
965 883
2 0 22 0 0 4096 0 69 0 0 118 2
279 104
279 59
2 1 2 0 0 0 0 25 67 0 0 5
313 179
279 179
279 138
238 138
238 147
3 0 22 0 0 12288 0 25 0 0 124 5
313 188
295 188
295 59
633 59
633 87
8 6 23 0 0 24704 0 78 25 0 0 8
753 935
771 935
771 1016
450 1016
450 901
32 901
32 215
313 215
9 0 24 0 0 4096 0 78 0 0 61 2
753 926
763 926
6 10 24 0 0 12416 0 78 78 0 0 6
687 926
668 926
668 949
763 949
763 917
753 917
7 5 25 0 0 8320 0 25 78 0 0 8
313 224
42 224
42 889
459 889
459 1006
659 1006
659 917
687 917
4 8 26 0 0 24704 0 78 25 0 0 8
687 908
649 908
649 996
468 996
468 877
54 877
54 233
313 233
13 9 11 0 0 24704 0 76 25 0 0 8
965 893
1026 893
1026 1053
410 1053
410 943
65 943
65 242
313 242
10 14 27 0 0 8320 0 25 76 0 0 8
313 251
76 251
76 932
419 932
419 1044
1018 1044
1018 903
965 903
15 11 28 0 0 24704 0 76 25 0 0 8
965 913
1009 913
1009 1035
430 1035
430 922
88 922
88 260
313 260
1 0 2 0 0 0 0 84 0 0 73 2
864 969
864 987
7 2 12 0 0 8320 0 76 84 0 0 3
902 913
864 913
864 933
6 0 3 0 0 0 0 77 0 0 77 4
540 913
514 913
514 839
619 839
4 5 16 0 0 0 0 77 77 0 0 4
540 895
532 895
532 904
540 904
1 0 2 0 0 0 0 6 0 0 75 2
604 1080
604 988
1 0 2 0 0 0 0 8 0 0 75 2
619 959
619 988
8 0 2 0 0 0 0 76 0 0 75 5
902 923
918 923
918 987
784 987
784 988
7 0 2 0 0 0 0 78 0 0 75 3
687 935
678 935
678 988
8 1 2 0 0 12288 0 77 7 0 0 5
540 931
526 931
526 988
784 988
784 922
2 0 3 0 0 0 0 7 0 0 77 2
784 904
784 881
16 14 3 0 0 0 0 77 78 0 0 7
606 868
606 867
619 867
619 839
784 839
784 881
753 881
1 2 29 0 0 0 0 78 78 0 0 4
687 881
675 881
675 890
687 890
3 1 4 0 0 0 0 78 76 0 0 6
687 899
664 899
664 852
891 852
891 853
902 853
9 1 30 0 0 8320 0 76 16 0 0 6
965 853
1027 853
1027 606
864 606
864 630
879 630
3 16 31 0 0 4224 0 17 25 0 0 4
684 697
131 697
131 305
313 305
3 17 32 0 0 8320 0 18 25 0 0 4
684 675
140 675
140 314
313 314
0 18 34 0 0 8320 0 0 25 84 0 5
822 647
822 790
151 790
151 323
313 323
2 1 34 0 0 0 0 15 85 0 0 6
879 647
822 647
822 658
823 658
823 622
742 622
3 19 35 0 0 12416 0 15 25 0 0 6
879 661
834 661
834 779
159 779
159 332
313 332
3 0 36 0 0 12416 0 1 0 0 95 4
878 683
869 683
869 768
566 768
2 0 15 0 0 0 0 9 0 0 92 4
956 712
982 712
982 713
997 713
5 1 37 0 0 4224 0 1 9 0 0 4
908 713
922 713
922 712
936 712
2 0 15 0 0 0 0 10 0 0 93 2
767 727
784 727
2 0 15 0 0 0 0 11 0 0 93 2
600 753
611 753
0 1 36 0 0 0 0 0 11 95 0 4
566 752
570 752
570 753
580 753
0 4 15 0 0 0 0 0 1 93 0 5
784 753
784 752
997 752
997 689
908 689
4 4 15 0 0 0 0 19 17 0 0 6
548 728
611 728
611 753
784 753
784 703
714 703
2 20 38 0 0 8320 0 19 25 0 0 4
518 708
171 708
171 341
313 341
3 5 36 0 0 0 0 19 19 0 0 6
518 722
502 722
502 768
566 768
566 752
548 752
1 1 2 0 0 0 0 12 15 0 0 5
848 688
848 676
847 676
847 654
879 654
1 0 2 0 0 0 0 17 0 0 98 2
684 690
652 690
1 1 2 0 0 0 0 13 18 0 0 3
652 707
652 668
684 668
1 1 2 0 0 0 0 14 19 0 0 3
473 735
473 715
518 715
12 0 2 0 0 0 0 21 0 0 107 3
445 599
486 599
486 651
21 7 43 0 0 8320 0 25 21 0 0 4
313 350
181 350
181 617
379 617
5 23 39 0 0 8320 0 21 25 0 0 4
379 599
199 599
199 368
313 368
22 6 44 0 0 8320 0 25 21 0 0 4
313 359
190 359
190 608
379 608
24 3 40 0 0 8320 0 25 21 0 0 4
313 377
209 377
209 581
379 581
2 25 45 0 0 8320 0 21 25 0 0 4
379 572
217 572
217 386
313 386
26 1 46 0 0 8320 0 25 21 0 0 4
313 395
227 395
227 563
379 563
1 0 2 0 0 0 0 75 0 0 109 3
532 596
532 651
307 651
2 16 3 0 0 0 0 75 21 0 0 4
532 578
533 578
533 563
445 563
1 8 2 0 0 0 0 74 21 0 0 3
307 657
307 626
379 626
1 0 2 0 0 0 0 73 0 0 129 3
753 584
753 592
734 592
0 2 22 0 0 0 0 0 73 124 0 3
745 488
753 488
753 566
1 0 2 0 0 0 0 72 0 0 128 3
649 465
649 469
624 469
0 2 22 0 0 0 0 0 72 125 0 3
633 366
649 366
649 447
1 0 2 0 0 0 0 71 0 0 127 3
763 315
763 322
734 322
2 0 22 0 0 0 0 71 0 0 123 3
763 297
763 217
745 217
2 0 22 0 0 0 0 70 0 0 124 2
651 164
651 87
0 1 2 0 0 0 0 0 70 126 0 3
621 191
651 191
651 182
1 0 22 0 0 0 0 68 0 0 58 3
238 105
238 59
295 59
0 1 2 0 0 0 0 0 34 122 0 3
984 227
984 73
1002 73
1 0 2 0 0 0 0 52 0 0 122 2
1000 358
984 358
1 0 2 0 0 0 0 61 0 0 122 2
1000 491
984 491
1 1 2 0 0 8320 0 43 66 0 0 5
1002 227
984 227
984 491
985 491
985 581
20 0 22 0 0 0 0 20 0 0 124 2
724 217
745 217
20 20 22 0 0 8192 0 24 22 0 0 4
612 87
745 87
745 488
725 488
20 0 22 0 0 0 0 23 0 0 124 4
617 367
617 366
633 366
633 87
11 0 2 0 0 0 0 24 0 0 195 4
612 168
621 168
621 191
532 191
11 1 2 0 0 0 0 20 28 0 0 4
724 298
734 298
734 322
650 322
1 11 2 0 0 0 0 27 23 0 0 4
533 469
625 469
625 448
617 448
1 11 2 0 0 0 0 26 22 0 0 4
648 592
734 592
734 569
725 569
2 10 67 0 0 4224 0 60 61 0 0 2
900 572
1000 572
2 9 68 0 0 12416 0 59 61 0 0 4
878 556
912 556
912 563
1000 563
2 8 69 0 0 12416 0 58 61 0 0 4
901 542
919 542
919 554
1000 554
2 7 70 0 0 12416 0 57 61 0 0 4
877 524
926 524
926 545
1000 545
2 6 71 0 0 12416 0 62 61 0 0 4
900 511
934 511
934 536
1000 536
2 5 72 0 0 4224 0 63 61 0 0 4
877 497
940 497
940 527
1000 527
2 4 73 0 0 12416 0 64 61 0 0 4
899 482
948 482
948 518
1000 518
1 12 74 0 0 12416 0 60 22 0 0 4
880 572
808 572
808 560
725 560
13 1 75 0 0 8320 0 22 59 0 0 5
725 551
725 550
844 550
844 556
858 556
1 14 76 0 0 4224 0 58 22 0 0 2
881 542
725 542
15 1 77 0 0 4224 0 22 57 0 0 4
725 533
843 533
843 524
857 524
3 2 78 0 0 12416 0 61 65 0 0 4
1000 509
956 509
956 466
877 466
16 1 79 0 0 4224 0 22 62 0 0 4
725 524
815 524
815 511
880 511
17 1 80 0 0 4224 0 22 63 0 0 4
725 515
801 515
801 497
857 497
18 1 81 0 0 12416 0 22 64 0 0 4
725 506
792 506
792 482
879 482
19 1 82 0 0 12416 0 22 65 0 0 4
725 497
783 497
783 466
857 466
2 10 83 0 0 4224 0 51 52 0 0 2
878 439
1000 439
2 9 84 0 0 12416 0 50 52 0 0 4
898 423
914 423
914 430
1000 430
2 8 85 0 0 12416 0 49 52 0 0 4
879 408
922 408
922 421
1000 421
2 7 86 0 0 12416 0 48 52 0 0 4
898 394
931 394
931 412
1000 412
2 6 87 0 0 4224 0 53 52 0 0 4
879 379
941 379
941 403
1000 403
2 5 88 0 0 4224 0 54 52 0 0 4
898 364
951 364
951 394
1000 394
2 4 89 0 0 4224 0 55 52 0 0 4
880 348
962 348
962 385
1000 385
1 12 90 0 0 4224 0 51 23 0 0 2
858 439
617 439
13 1 91 0 0 4224 0 23 50 0 0 4
617 430
835 430
835 423
878 423
1 14 92 0 0 12416 0 49 23 0 0 4
859 408
827 408
827 421
617 421
15 1 93 0 0 4224 0 23 48 0 0 4
617 412
817 412
817 394
878 394
3 2 94 0 0 12416 0 52 56 0 0 4
1000 376
972 376
972 331
898 331
16 1 95 0 0 4224 0 23 53 0 0 4
617 403
807 403
807 379
859 379
17 1 96 0 0 4224 0 23 54 0 0 4
617 394
798 394
798 364
878 364
18 1 97 0 0 4224 0 23 55 0 0 4
617 385
789 385
789 348
860 348
19 1 98 0 0 4224 0 23 56 0 0 4
617 376
777 376
777 331
878 331
2 10 99 0 0 4224 0 42 43 0 0 2
879 308
1002 308
2 9 100 0 0 12416 0 41 43 0 0 4
899 293
911 293
911 299
1002 299
2 8 101 0 0 12416 0 40 43 0 0 4
879 277
918 277
918 290
1002 290
2 7 102 0 0 12416 0 39 43 0 0 4
899 261
926 261
926 281
1002 281
2 6 103 0 0 12416 0 44 43 0 0 4
881 244
935 244
935 272
1002 272
2 5 104 0 0 12416 0 45 43 0 0 4
898 228
944 228
944 263
1002 263
2 4 105 0 0 4224 0 46 43 0 0 4
880 212
953 212
953 254
1002 254
1 12 106 0 0 12416 0 42 20 0 0 4
859 308
798 308
798 289
724 289
13 1 107 0 0 4224 0 20 41 0 0 4
724 280
807 280
807 293
879 293
1 14 108 0 0 12416 0 40 20 0 0 4
859 277
817 277
817 271
724 271
15 1 109 0 0 4224 0 20 39 0 0 4
724 262
864 262
864 261
879 261
3 2 110 0 0 12416 0 43 47 0 0 4
1002 245
963 245
963 196
898 196
16 1 111 0 0 4224 0 20 44 0 0 4
724 253
817 253
817 244
861 244
17 1 112 0 0 4224 0 20 45 0 0 4
724 244
808 244
808 228
878 228
18 1 113 0 0 4224 0 20 46 0 0 4
724 235
798 235
798 212
860 212
19 1 114 0 0 12416 0 20 47 0 0 4
724 226
786 226
786 196
878 196
2 10 115 0 0 4224 0 35 34 0 0 4
879 179
959 179
959 154
1002 154
2 9 116 0 0 12416 0 36 34 0 0 4
899 164
947 164
947 145
1002 145
2 8 117 0 0 12416 0 37 34 0 0 4
882 149
936 149
936 136
1002 136
2 7 118 0 0 12416 0 38 34 0 0 4
902 132
922 132
922 127
1002 127
2 6 119 0 0 4224 0 33 34 0 0 2
882 118
1002 118
2 5 120 0 0 12416 0 32 34 0 0 4
903 103
923 103
923 109
1002 109
2 4 121 0 0 12416 0 31 34 0 0 4
883 87
935 87
935 100
1002 100
1 12 122 0 0 12416 0 35 24 0 0 4
859 179
775 179
775 159
612 159
13 1 123 0 0 4224 0 24 36 0 0 4
612 150
784 150
784 164
879 164
1 14 124 0 0 12416 0 37 24 0 0 4
862 149
796 149
796 141
612 141
15 1 125 0 0 4224 0 24 38 0 0 2
612 132
882 132
3 2 126 0 0 4224 0 34 30 0 0 4
1002 91
946 91
946 71
903 71
16 1 127 0 0 4224 0 24 33 0 0 4
612 123
793 123
793 118
862 118
17 1 128 0 0 4224 0 24 32 0 0 4
612 114
784 114
784 103
883 103
18 1 129 0 0 4224 0 24 31 0 0 4
612 105
773 105
773 87
863 87
19 1 130 0 0 4224 0 24 30 0 0 4
612 96
761 96
761 71
883 71
10 0 2 0 0 0 0 24 0 0 195 2
546 168
532 168
9 1 2 0 0 0 0 24 29 0 0 5
546 159
532 159
532 191
533 191
533 194
10 0 2 0 0 0 0 20 0 0 197 2
658 298
651 298
9 1 2 0 0 0 0 20 28 0 0 5
658 289
651 289
651 298
650 298
650 322
10 0 2 0 0 0 0 23 0 0 199 2
551 448
533 448
9 1 2 0 0 0 0 23 27 0 0 3
551 439
533 439
533 469
10 0 2 0 0 0 0 22 0 0 201 2
659 569
648 569
1 9 2 0 0 0 0 26 22 0 0 3
648 592
648 560
659 560
8 41 139 0 0 12416 0 23 25 0 0 4
551 430
468 430
468 377
379 377
42 7 140 0 0 4224 0 25 23 0 0 4
379 368
477 368
477 421
551 421
6 43 141 0 0 12416 0 23 25 0 0 4
551 412
488 412
488 359
379 359
44 5 142 0 0 4224 0 25 23 0 0 4
379 350
498 350
498 403
551 403
4 45 143 0 0 12416 0 23 25 0 0 4
551 394
506 394
506 341
379 341
46 3 144 0 0 4224 0 25 23 0 0 4
379 332
516 332
516 385
551 385
2 47 145 0 0 12416 0 23 25 0 0 4
551 376
525 376
525 323
379 323
48 1 146 0 0 4224 0 25 23 0 0 4
379 314
534 314
534 367
551 367
8 49 147 0 0 12416 0 20 25 0 0 4
658 280
617 280
617 305
379 305
50 7 148 0 0 4224 0 25 20 0 0 4
379 296
607 296
607 271
658 271
6 51 149 0 0 12416 0 20 25 0 0 4
658 262
596 262
596 287
379 287
52 5 150 0 0 4224 0 25 20 0 0 4
379 278
585 278
585 253
658 253
4 53 151 0 0 12416 0 20 25 0 0 4
658 244
575 244
575 269
379 269
54 3 152 0 0 4224 0 25 20 0 0 4
379 260
563 260
563 235
658 235
2 55 153 0 0 12416 0 20 25 0 0 4
658 226
551 226
551 251
379 251
56 1 154 0 0 4224 0 25 20 0 0 4
379 242
540 242
540 217
658 217
8 57 155 0 0 12416 0 24 25 0 0 4
546 150
515 150
515 233
379 233
58 7 156 0 0 4224 0 25 24 0 0 4
379 224
504 224
504 141
546 141
6 59 157 0 0 12416 0 24 25 0 0 4
546 132
494 132
494 215
379 215
60 5 158 0 0 4224 0 25 24 0 0 4
379 206
484 206
484 123
546 123
4 61 159 0 0 12416 0 24 25 0 0 4
546 114
475 114
475 197
379 197
62 3 160 0 0 4224 0 25 24 0 0 4
379 188
465 188
465 105
546 105
2 63 161 0 0 4224 0 24 25 0 0 4
546 96
455 96
455 179
379 179
64 1 162 0 0 12416 0 25 24 0 0 4
379 170
443 170
443 87
546 87
62
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 15
674 601 786 624
679 605 784 620
15 POWER ON ENABLE
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 16
339 522 458 545
344 526 456 541
16 E.STOP LED DRIVE
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 18
327 513 460 536
332 517 458 532
18 POWER ON LED DRIVE
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 18
405 1217 538 1240
410 1221 536 1236
18 POWER ON SENSE-OUT
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 18
616 1230 749 1253
621 1233 747 1248
18 E.STOP PILOT LIGHT
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 17
119 984 231 1007
126 989 232 1004
17 POWER ON SENSE-IN
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 23
84 195 252 218
89 199 250 214
23 CAMERA LIGHT ON/OFF-OUT
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 22
85 186 246 209
90 190 244 205
22 CAMERA LIGHT ON/OFF-IN
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
124 258 152 281
129 262 150 277
3 EN3
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
123 267 151 290
128 271 149 286
3 EN2
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
123 276 151 299
128 280 149 295
3 EN1
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
123 285 151 308
128 289 149 304
3 EN0
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 15
125 249 237 272
130 253 235 268
15 TOWER LIGHT RED
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 15
125 240 237 263
130 244 235 259
15 TOWER LIGHT YLW
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 15
127 231 239 254
132 235 237 250
15 TOWER LIGHT GRN
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 8
311 46 374 69
316 50 372 65
8 VCC(+5V)
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 4
394 158 429 181
399 162 427 177
4 Z1-A
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
394 168 436 191
399 172 434 187
5 Z1-*A
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 4
395 176 430 199
400 180 428 195
4 ZI-B
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
393 186 435 209
398 190 433 205
5 Z1-*B
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 4
395 195 430 218
400 199 428 214
4 T1-A
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
395 204 437 227
400 208 435 223
5 T1-*A
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 4
396 213 431 236
401 217 429 232
4 T1-B
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
394 221 436 244
399 225 434 240
5 T1-*B
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 4
396 230 431 253
401 234 429 249
4 Z2-A
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
396 239 438 262
401 243 436 258
5 Z2-*A
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 4
396 248 431 271
401 252 429 267
4 Z2-B
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
396 257 438 280
401 261 436 276
5 Z2-*B
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 4
396 266 431 289
401 270 429 285
4 T2-A
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
395 275 437 298
400 279 435 294
5 T2-*A
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 4
396 284 431 307
401 288 429 303
4 T2-B
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
395 293 437 316
400 297 435 312
5 T2-*B
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 4
395 303 430 326
400 307 428 322
4 XR-A
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
395 312 437 335
400 316 435 331
5 XR-*A
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 4
397 321 432 344
402 325 430 340
4 XR-B
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
396 329 438 352
401 333 436 348
5 XR-*B
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 4
398 338 433 361
403 342 431 357
4 YR-A
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
397 348 439 371
402 352 437 367
5 YR-*A
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 4
397 357 432 380
402 361 430 376
4 YR-B
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
396 366 438 389
401 370 436 385
5 YR-*B
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
395 375 423 398
400 379 421 394
3 X-H
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 4
396 383 431 406
401 387 429 402
4 X-*H
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
384 410 412 433
389 414 410 429
3 Y-H
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 4
379 420 414 443
384 424 412 439
4 Y-*H
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 4
264 384 299 407
269 388 297 403
4 Z1-H
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
263 375 305 398
268 379 303 394
5 Z1-*H
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 4
265 348 300 371
270 352 298 367
4 Z2-H
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
263 340 305 363
268 344 303 359
5 Z2-*H
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
396 392 417 415
401 396 415 411
2 XH
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
397 402 418 425
402 406 416 421
2 YH
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
265 368 293 391
270 372 291 387
3 Z1H
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
265 357 293 380
270 361 291 376
3 Z2H
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 9
198 329 260 352
204 334 260 349
9 E.STOP SW
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 8
200 320 256 343
206 325 256 340
8 RESET SW
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 12
200 311 281 334
206 316 281 331
12 E.STOP SENSE
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 12
863 593 944 616
869 598 944 613
12 P. ON ENABLE
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 17
138 293 250 316
144 298 250 313
17 AC SERVO POWER ON
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 20
136 303 267 326
143 308 268 323
20 Z1,Z2,T1,T2 POWER ON
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 8
126 213 189 236
131 217 187 232
8 DOOR SW1
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 8
126 222 189 245
131 226 187 241
8 DOOR SW2
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 10
126 204 203 227
131 208 201 223
10 DOOR SW OK
-11 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 4
262 429 297 452
267 433 295 448
4 +24V
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
