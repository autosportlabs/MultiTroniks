CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
20 130 30 100 9
0 66 800 572
7 5.000 V
7 5.000 V
3 GND
1000 10
24 100 0 1 1
20 Package,Description,
61 C:\PROGRAM FILES\MICROCODE ENGINEERING\CIRCUITMAKER 6\BOM.DAT
0 7
0 66 800 572
12058642 80
2
38 AC SERVOPACK INTERFACE CIRCUIT DIAGRAM
50 MULTITRONIKS
ONE FREDERICK ROAD, WARREN, NJ 07059
0
0
4 LVX2
12
10 Polar Cap~
219 268 471 0 2 5
0 3 2
0
0 0 832 180
5 100uF
-22 -18 13 -10
2 C1
-11 -28 3 -20
0
0
11 %D %1 %2 %V
0
0
7 RB.2/.4
5

0 1 2 1 2 -1610612675
67 0 0 0 1 0 0 0
1 C
8953 0 0
0
0
7 Ground~
168 216 491 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4441 0 0
0
0
5 CON20
94 556 410 0 20 41
0 2 23 21 2 19 17 7 5 2
3 24 22 2 20 18 2 6 4 2
3
5 CON20
1 0 4736 0
4 CONN
-14 -66 14 -58
2 J3
-7 -66 7 -58
0
0
0
0
0
5 IDC20
41

0 1 3 5 7 9 11 13 15 17
19 2 4 6 8 10 12 14 16 18
20 1 3 5 7 9 11 13 15 17
19 2 4 6 8 10 12 14 16 18
20 0
0 0 0 0 1 0 0 0
1 J
3618 0 0
0
0
7 Ground~
168 572 211 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6153 0 0
0
0
7 Ground~
168 483 513 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5394 0 0
0
0
7 Ground~
168 403 263 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7734 0 0
0
0
7 Ground~
168 110 174 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9914 0 0
0
0
7 Ground~
168 110 431 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3747 0 0
0
0
4 2003
94 359 221 0 16 33
0 15 62 63 64 65 66 14 2 12
67 68 69 70 71 11 3
4 2003
2 0 6528 512
2 U1
-8 -55 6 -47
2 U1
-8 -65 6 -57
0
0
0
0
0
5 DIP16
33

0 1 2 3 4 5 6 7 8 16
15 14 13 12 11 10 9 1 2 3
4 5 6 7 8 16 15 14 13 12
11 10 9 0
0 0 0 512 1 1 0 0
1 A
3549 0 0
0
0
5 CON12
94 102 145 0 12 25
0 24 23 22 21 13 9 2 11 3
7 6 72
5 CON12
3 0 4480 0
2 J1
-36 -109 -22 -101
2 J1
-31 -120 -17 -112
0
0
0
0
0
7 MOLEX12
25

0 1 2 3 4 5 6 7 8 9
10 11 12 1 2 3 4 5 6 7
8 9 10 11 12 0
0 0 0 512 1 1 0 0
1 J
7931 0 0
0
0
5 CON10
94 626 193 0 10 21
0 13 14 16 15 73 2 9 2 8
74
5 CON10
4 0 4480 0
2 J4
-17 -60 -3 -52
2 J4
-17 -70 -3 -62
0
0
0
0
0
5 IDC10
21

0 2 4 6 8 10 1 3 5 7
9 2 4 6 8 10 1 3 5 7
9 0
0 0 0 512 1 0 0 0
1 A
9325 0 0
0
0
5 CON12
94 100 405 0 12 25
0 20 19 18 17 16 8 2 12 3
5 4 75
5 CON12
5 0 12928 0
5 CON12
-41 -110 -6 -102
2 J2
-39 -114 -25 -106
0
0
0
0
0
7 MOLEX12
25

0 1 2 3 4 5 6 7 8 9
10 11 12 1 2 3 4 5 6 7
8 9 10 11 12 0
0 0 0 512 1 0 0 0
1 J
8903 0 0
0
0
38
1 0 3 0 0 4096 0 1 0 0 5 2
275 471
302 471
2 1 2 0 0 4096 0 1 2 0 0 3
258 471
216 471
216 485
0 0 2 0 0 12416 0 0 0 7 14 4
632 444
631 444
631 492
483 492
20 0 3 0 0 12288 0 3 0 0 5 4
578 454
611 454
611 471
509 471
0 10 3 0 0 8192 0 0 3 21 0 5
302 395
302 471
509 471
509 454
534 454
9 0 2 0 0 0 0 3 0 0 14 2
534 444
483 444
19 0 2 0 0 0 0 3 0 0 12 3
578 444
632 444
632 414
11 18 4 0 0 12416 0 12 3 0 0 6
93 415
321 415
321 482
621 482
621 434
578 434
10 8 5 0 0 4224 0 12 3 0 0 4
93 405
339 405
339 434
534 434
11 17 6 0 0 12416 0 10 3 0 0 6
95 155
200 155
200 325
653 325
653 424
578 424
10 7 7 0 0 20608 0 10 3 0 0 6
95 145
212 145
212 260
231 260
231 424
534 424
16 13 2 0 0 0 0 3 3 0 0 4
578 414
632 414
632 384
578 384
4 0 2 0 0 0 0 3 0 0 14 2
534 394
483 394
1 1 2 0 0 0 0 3 5 0 0 3
534 364
483 364
483 507
8 0 2 0 0 0 0 11 0 0 16 2
584 174
572 174
6 1 2 0 0 0 0 11 4 0 0 3
584 153
572 153
572 205
6 9 8 0 0 12416 0 12 11 0 0 6
93 365
108 365
108 276
429 276
429 183
584 183
6 7 9 0 0 12416 0 10 11 0 0 4
95 105
327 105
327 163
584 163
0 0 10 0 0 4224 0 0 0 0 0 3
599 67
599 66
598 66
8 15 11 0 0 4224 0 10 9 0 0 4
95 125
224 125
224 245
326 245
0 9 3 0 0 8320 0 0 12 22 0 3
302 255
302 395
93 395
9 16 3 0 0 0 0 10 9 0 0 4
95 135
302 135
302 255
326 255
8 9 12 0 0 12416 0 12 9 0 0 4
93 385
99 385
99 185
326 185
1 5 13 0 0 12416 0 11 10 0 0 4
649 153
652 153
652 95
95 95
7 2 14 0 0 12416 0 9 11 0 0 6
389 245
400 245
400 125
662 125
662 163
649 163
4 1 15 0 0 12416 0 11 9 0 0 6
649 183
653 183
653 234
411 234
411 185
389 185
3 5 16 0 0 20608 0 11 12 0 0 6
649 173
662 173
662 255
441 255
441 355
93 355
4 6 17 0 0 12416 0 12 3 0 0 6
93 345
118 345
118 384
355 384
355 414
534 414
3 15 18 0 0 4224 0 12 3 0 0 4
93 335
642 335
642 404
578 404
2 5 19 0 0 12416 0 12 3 0 0 6
93 325
145 325
145 374
370 374
370 404
534 404
7 1 2 0 0 0 0 12 8 0 0 3
93 375
110 375
110 425
14 1 20 0 0 12416 0 3 12 0 0 6
578 394
618 394
618 345
157 345
157 315
93 315
4 3 21 0 0 8320 0 10 3 0 0 6
95 85
243 85
243 316
385 316
385 384
534 384
12 3 22 0 0 12416 0 3 10 0 0 6
578 374
608 374
608 306
252 306
252 75
95 75
2 2 23 0 0 8320 0 10 3 0 0 6
95 65
261 65
261 297
399 297
399 374
534 374
1 11 24 0 0 12416 0 10 3 0 0 6
95 55
272 55
272 287
600 287
600 364
578 364
8 1 2 0 0 0 0 9 6 0 0 3
389 255
403 255
403 257
7 1 2 0 0 0 0 10 7 0 0 3
95 115
110 115
110 168
56
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 5
660 153 689 168
664 157 688 168
5 X INH
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 6
659 164 695 179
663 168 694 179
6 Y REF+
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 5
660 174 689 189
664 178 688 189
5 Y INH
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 3
559 139 585 154
563 143 584 154
3 GND
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 3
547 162 573 177
551 166 572 177
3 GND
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 6
516 149 551 164
520 153 550 164
6 X REF-
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 6
516 169 551 184
520 173 550 184
6 Y REF-
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 3
492 351 518 366
496 355 517 366
3 GND
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 2
579 351 597 366
583 354 596 365
2 XA
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 3
496 360 517 375
500 364 516 375
3 *XA
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 6
7 46 45 61
11 50 44 61
6 22 PBO
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 7
7 57 48 72
11 61 47 72
7 23 *PBO
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 6
6 67 44 82
10 71 43 82
6 20 PAO
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 7
7 77 48 92
11 81 47 92
7 21 *PAO
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 7
7 87 47 102
11 91 46 102
7 1 T-REF
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 4
7 97 32 112
11 101 31 112
4 2 SG
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 5
6 107 36 122
10 111 35 122
5 19 SG
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 7
6 116 46 131
10 120 45 131
7 14 S-ON
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 6
14 306 52 321
18 310 51 321
6 35 PBO
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 7
13 316 54 331
17 320 53 331
7 36 *PBO
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 6
14 326 52 341
18 330 51 341
6 33 PAO
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 7
14 338 55 353
18 342 54 353
7 34 *PAO
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 7
13 347 53 362
17 351 52 362
7 9 T-REF
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 5
13 357 43 372
17 361 42 372
5 10 SG
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 4
13 367 38 382
17 371 37 382
4 1 SG
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 7
12 377 52 392
16 381 51 392
7 40 S-ON
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 10
12 387 60 402
16 390 59 401
10 47 +24V IN
-13 0 0 0 400 0 0 0 0 3 2 1 18
15 Times New Roman
0 0 0 44
655 350 750 425
659 354 749 414
44 TO MOTION
CONTROLLER
INTERFACE
BOARD  J13
-13 0 0 0 400 0 0 0 0 3 2 1 18
15 Times New Roman
0 0 0 30
707 136 793 193
711 140 792 185
30 TO I/O
INTERFACE 
BOARD  J11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
7 269 31 293
11 273 27 289
2 TO
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
44 10 68 34
48 14 64 30
2 TO
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 10
6 127 54 142
10 131 53 142
10 13 +24V IN
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
32 269 216 293
36 273 212 289
22 Y AXIS 1CN(SGDB-15ADG)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
66 9 242 33
70 13 238 29
21 X AXIS 1CN(SGDA-04AS)
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 6
660 143 696 158
664 147 695 158
6 X REF+
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 3
499 401 520 416
503 405 519 416
3 *YB
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 2
581 391 599 406
585 395 598 406
2 YB
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 3
498 391 519 406
502 395 518 406
3 *YA
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 2
581 382 599 397
585 386 598 397
2 YA
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 3
496 381 522 396
500 385 521 396
3 GND
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 3
577 371 603 386
581 375 602 386
3 GND
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 3
496 371 517 386
500 375 516 386
3 *XB
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 2
579 362 597 377
583 366 596 377
2 XB
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 6
7 137 45 152
11 141 44 152
6 24 PCO
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 7
7 146 48 161
11 150 47 161
7 25 *PCO
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 6
13 396 51 411
17 400 50 411
6 19 PCO
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 7
13 406 54 421
17 410 53 421
7 20 *PCO
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 3
580 403 606 418
584 406 605 417
3 GND
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 6
493 411 529 426
497 415 528 426
6   XPCO
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 5
577 411 612 426
581 415 611 426
5 *XPCO
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 4
495 421 527 436
499 425 526 436
4 YPCO
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 5
579 421 614 436
583 425 613 436
5 *YPCO
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 3
499 431 525 446
503 435 524 446
3 GND
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 3
584 431 610 446
588 435 609 446
3 GND
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 4
584 441 609 456
588 445 608 456
4 +24V
-9 0 0 0 400 0 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 4
500 441 525 456
504 445 524 456
4 +24V
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
