CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 40 9
20 78 780 559
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
61 C:\PROGRAM FILES\MICROCODE ENGINEERING\CIRCUITMAKER 6\BOM.DAT
0 7
20 78 780 559
146276370 80
2
31 Title:KEY BOARD EXTENSION CACLE
51 MULTITRONIKS
ONE FREDERICK ROAD - WARREN, NJ 07059
10 09-17-1998
0
4 LVX2
2
4 PLUG
94 803 306 0 1 3
0 0
4 PLUG
1 0 0 0
0
2 U1
-7 -29 7 -21
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
1 P
8953 0 0
0
0
7 SOCKET~
94 108 305 0 6 13
0 2 2 2 2 2 2
7 SOCKET~
2 0 2560 0
0
2 U2
-6 -57 8 -49
0
0
0
0
0
0
13

0 3 5 2 4 1 -195123 3 5 2
4 1 -195123 0
0 0 0 0 1 1 0 0
1 C
4441 0 0
0
0
7
0 6 2 0 0 12288 0 0 2 2 0 6
227 305
225 305
225 240
63 240
63 307
81 307
0 1 2 0 0 0 0 0 2 3 0 5
227 306
227 305
219 305
219 279
108 279
0 2 2 0 0 0 0 0 2 4 0 4
227 306
215 306
215 292
128 292
0 5 2 0 0 0 0 0 2 5 0 5
227 307
227 306
219 306
219 334
108 334
0 4 2 0 0 0 0 0 2 6 0 5
227 306
227 307
214 307
214 321
127 321
0 3 2 0 0 0 0 0 2 7 0 2
228 306
135 306
0 0 2 0 0 12416 0 0 0 0 0 4
712 302
228 302
228 310
713 310
11
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
151 322 201 343
155 326 197 341
5 BROWN
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
164 295 197 316
167 299 192 314
3 RED
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
146 268 204 289
150 272 200 287
6 ORANGE
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
148 310 206 331
152 313 202 328
6 YELLOW
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
153 281 203 302
157 284 199 299
5 GREEN
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
150 230 200 251
154 233 196 248
5 BLACK
-16 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 15
861 358 1008 386
865 362 1003 380
15 PIN ASSIGHNMENT
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 64
860 385 960 496
864 388 956 478
64   1.BROWN
  2.RED
  3.ORANGE
  4.YELLOW
  5.GREEN
GND.BLACK
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 13
757 253 873 292
761 256 869 286
13 PLUG P#18665-
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 33
381 266 539 305
385 270 535 300
33 CABLE P#19274-
LENGTH 120 INCHES
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 15
60 360 193 381
63 364 188 379
15 SOCKET P#18666-
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
