CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 60 30 100 9
0 68 800 600
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
65 C:\PROGRAM FILES\MICROCODE ENGINEERING\CIRCUITMAKER 6 PRO\BOM.DAT
0 7
0 68 800 600
144179218 0
0
6 Title:
5 Name:
0
0
0
19
6 Diode~
219 561 203 0 2 5
0 4 3
0
0 0 848 90
5 DIODE
11 0 46 8
2 D1
22 -10 36 -2
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
8953 0 0
0
0
14 NO PushButton~
191 99 319 0 2 5
0 13 3
0
0 0 4720 0
0
2 S1
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
4441 0 0
0
0
5 SIP2~
219 634 192 0 2 5
0 3 4
0
0 0 624 0
4 CONN
9 2 37 10
2 J2
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 -1610612472
0 0 0 0 1 0 0 0
1 J
3618 0 0
0
0
5 SIP3~
219 113 249 0 3 7
0 2 6 3
0
0 0 624 180
4 CONN
-13 -25 15 -17
2 J1
-10 -26 4 -18
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 -1610612488
0 0 0 0 1 0 0 0
1 J
6153 0 0
0
0
12 NPN Trans:C~
219 408 347 0 3 7
0 7 9 2
0
0 0 848 0
6 2N3904
10 7 52 15
2 Q5
15 -4 29 4
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 0 0 0
1 Q
5394 0 0
0
0
12 NPN Trans:C~
219 504 307 0 3 7
0 4 7 2
0
0 0 848 0
6 2N3904
10 9 52 17
2 Q2
16 -3 30 5
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 0 0 0
1 Q
7734 0 0
0
0
12 PNP Trans:C~
219 504 227 0 3 7
0 4 12 3
0
0 0 848 692
6 2N3906
11 7 53 15
2 Q1
16 -5 30 3
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
113 0 0 0 1 0 0 0
1 Q
9914 0 0
0
0
12 NPN Trans:C~
219 226 327 0 3 7
0 8 5 2
0
0 0 976 0
6 2N3904
7 23 49 31
2 Q4
15 -3 29 5
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -1610612700
81 0 0 0 1 0 0 0
1 Q
3747 0 0
0
0
12 NPN Trans:C~
219 337 291 0 3 7
0 11 10 2
0
0 0 848 0
6 2N3904
10 9 52 17
2 Q3
16 -3 30 5
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -1610612596
81 0 0 0 1 0 0 0
1 Q
3549 0 0
0
0
7 Ground~
168 413 404 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7931 0 0
0
0
9 Resistor~
219 183 367 0 3 5
0 2 5 -1
0
0 0 880 90
3 18k
5 0 26 8
2 R7
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612676
82 0 0 0 1 0 0 0
1 R
9325 0 0
0
0
9 Resistor~
219 161 247 0 2 5
0 6 5
0
0 0 880 0
4 5.6k
-14 -14 14 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612676
82 0 0 0 1 0 0 0
1 R
8903 0 0
0
0
9 Resistor~
219 413 264 0 2 5
0 7 3
0
0 0 880 90
4 5.6k
4 0 32 8
3 R10
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612720
82 0 0 0 1 0 0 0
1 R
3834 0 0
0
0
9 Resistor~
219 297 347 0 2 5
0 8 9
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R9
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612676
82 0 0 0 1 0 0 0
1 R
3363 0 0
0
0
9 Resistor~
219 291 291 0 2 5
0 8 10
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612596
82 0 0 0 1 0 0 0
1 R
7668 0 0
0
0
9 Resistor~
219 231 207 0 2 5
0 8 3
0
0 0 880 90
3 18k
5 0 26 8
2 R6
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612696
82 0 0 0 1 0 0 0
1 R
4718 0 0
0
0
9 Resistor~
219 442 227 0 2 5
0 11 12
0
0 0 880 0
4 5.6k
-14 -14 14 -6
2 R5
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612720
82 0 0 0 1 0 0 0
1 R
3874 0 0
0
0
9 Resistor~
219 165 327 0 2 5
0 13 5
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612700
82 0 0 0 1 0 0 0
1 R
6671 0 0
0
0
9 Resistor~
219 342 182 0 2 5
0 11 3
0
0 0 880 90
4 5.6k
1 0 29 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612720
82 0 0 0 1 0 0 0
1 R
3789 0 0
0
0
31
1 0 4 0 0 0 0 1 0 0 28 2
561 213
561 267
2 0 3 0 0 4096 0 1 0 0 10 2
561 193
561 149
1 0 2 0 0 0 0 11 0 0 5 3
183 385
183 398
184 398
2 0 5 0 0 4096 0 11 0 0 29 2
183 349
183 327
1 0 2 0 0 8320 0 4 0 0 22 4
120 256
134 256
134 398
233 398
2 0 3 0 0 8192 0 2 0 0 7 4
82 327
65 327
65 149
134 149
3 0 3 0 0 0 0 4 0 0 23 4
120 238
134 238
134 149
231 149
2 0 5 0 0 8320 0 12 0 0 29 3
179 247
208 247
208 327
2 1 6 0 0 4224 0 4 12 0 0 2
120 247
143 247
1 0 3 0 0 0 0 3 0 0 23 4
622 188
617 188
617 149
509 149
2 0 3 0 0 0 0 13 0 0 23 2
413 246
413 149
1 0 2 0 0 0 0 10 0 0 16 2
413 398
413 398
2 0 3 0 0 0 0 19 0 0 23 2
342 164
342 149
2 0 7 0 0 4224 0 6 0 0 15 2
486 307
413 307
1 1 7 0 0 0 0 13 5 0 0 2
413 282
413 329
3 0 2 0 0 0 0 5 0 0 22 3
413 365
413 398
342 398
0 1 8 0 0 4096 0 0 14 20 0 3
273 291
273 347
279 347
2 2 9 0 0 4224 0 14 5 0 0 2
315 347
390 347
2 2 10 0 0 4224 0 15 9 0 0 2
309 291
319 291
0 1 8 0 0 0 0 0 15 24 0 2
231 291
273 291
1 0 11 0 0 4224 0 17 0 0 30 2
424 227
342 227
3 3 2 0 0 0 0 9 8 0 0 4
342 309
342 398
231 398
231 345
3 2 3 0 0 8320 0 7 16 0 0 4
509 209
509 149
231 149
231 189
1 1 8 0 0 4224 0 16 8 0 0 2
231 225
231 309
2 2 12 0 0 4224 0 17 7 0 0 2
460 227
486 227
3 0 2 0 0 0 0 6 0 0 16 3
509 325
509 398
413 398
1 0 4 0 0 0 0 6 0 0 28 2
509 289
509 267
1 2 4 0 0 128 0 7 3 0 0 5
509 245
509 267
617 267
617 197
622 197
2 2 5 0 0 0 0 18 8 0 0 2
183 327
208 327
1 1 11 0 0 0 0 9 19 0 0 2
342 273
342 200
1 1 13 0 0 4224 0 2 18 0 0 2
116 327
147 327
0
0
1 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
2316 1079360 100 100 0 0
0 0 0 0
299 97 460 167
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12401 0
4 10 1000
1
561 196
0 3 0 0 2	1 0 0 0
2820 8419392 100 100 0 0
77 66 767 186
0 334 800 600
767 66
77 66
767 66
767 186
0 0
0 0 0 0 0 0
12385 0
4 1e-006 50
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
