CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
650 290 30 120 9
0 66 796 576
7 5.000 V
7 5.000 V
3 GND
1000 10
24 100 0 1 0
20 Package,Description,
61 C:\PROGRAM FILES\MICROCODE ENGINEERING\CIRCUITMAKER 6\BOM.DAT
0 7
0 66 796 576
144179218 0
0
0
0
0
0
0
88
6 Diode~
219 641 990 0 2 5
0 19 20
0
0 0 64 90
5 DIODE
11 -5 46 3
2 D1
21 -15 35 -7
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
8953 0 0
0
0
6 Diode~
219 641 907 0 2 5
0 21 18
0
0 0 64 90
5 DIODE
11 -5 46 3
2 D2
21 -15 35 -7
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
4441 0 0
0
0
6 Diode~
219 641 831 0 2 5
0 22 17
0
0 0 64 90
5 DIODE
11 -5 46 3
2 D3
21 -15 35 -7
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3618 0 0
0
0
9 Rly sock~
94 651 907 0 16 33
0 78 79 2 2 21 80 81 18 82
83 84 85 86 87 88 89
8 Rly sock
1 0 0 0
0
0
0
0
0
0
0
0
33

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0
0 0 0 512 1 0 0 0
0
6153 0 0
0
0
9 Rly sock~
94 651 991 0 16 33
0 2 90 91 92 19 93 94 20 95
96 97 98 99 100 101 102
8 Rly sock
2 0 0 0
0
0
0
0
0
0
0
0
33

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0
0 0 0 512 1 0 0 0
0
5394 0 0
0
0
9 Rly sock~
94 651 829 0 16 33
0 103 104 2 2 22 105 106 17 107
108 109 110 111 112 113 114
8 Rly sock
3 0 0 0
0
0
0
0
0
0
0
0
33

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0
0 0 0 512 1 0 0 0
0
7734 0 0
0
0
6 Diode~
219 348 819 0 2 5
0 23 24
0
0 0 64 0
5 DIODE
-18 -18 17 -10
2 D4
-8 -28 6 -20
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 1 2 1 2 -1610612676
68 0 0 0 1 0 0 0
1 D
9914 0 0
0
0
5 Ter1~
94 1200 1165 0 1 3
0 28
4 Ter1
4 0 0 0
0
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3747 0 0
0
0
5 Ter1~
94 1200 1155 0 1 3
0 26
4 Ter1
5 0 0 0
0
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3549 0 0
0
0
5 Ter1~
94 1200 1145 0 1 3
0 11
4 Ter1
6 0 0 0
0
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
7931 0 0
0
0
5 Ter1~
94 1200 1137 0 1 3
0 12
4 Ter1
7 0 0 0
0
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
9325 0 0
0
0
5 Ter1~
94 1200 1127 0 1 3
0 13
4 Ter1
8 0 0 0
0
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
8903 0 0
0
0
5 Ter1~
94 1340 1202 0 1 3
0 27
4 Ter1
9 0 0 0
0
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3834 0 0
0
0
5 Ter1~
94 1340 1192 0 1 3
0 25
4 Ter1
10 0 0 0
0
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3363 0 0
0
0
5 Ter1~
94 1340 1182 0 1 3
0 14
4 Ter1
11 0 0 0
0
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
7668 0 0
0
0
5 Ter1~
94 1340 1172 0 1 3
0 15
4 Ter1
12 0 0 0
0
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
4718 0 0
0
0
5 Ter1~
94 1340 1162 0 1 3
0 16
4 Ter1
13 0 0 0
0
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3874 0 0
0
0
13 Relay Coil:C~
210 347 781 0 10 11
0 23 24 0 0 0 0 0 0 0
1
0
0 0 4192 0
7 24VCOIL
-24 10 25 18
2 X5
-7 -30 7 -22
0
0
24 *p=1 r=1
%D %1 %2 %I %S
0
11 alias:XCOIL
4 SIP2
5

0 1 2 1 2 0
88 0 0 0 1 0 0 0
3 RLY
6671 0 0
0
0
5 SIP2~
219 159 735 0 2 5
0 31 32
0
0 0 96 180
4 CONN
9 2 37 10
0
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 -1610612720
0 0 0 0 1 0 0 0
1 J
3789 0 0
0
0
10 TER BLOCK~
94 1232 243 0 2 5
0 115 116
10 TER BLOCK~
14 0 0 90
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
4871 0 0
0
0
10 TER BLOCK~
94 1243 243 0 2 5
0 117 118
10 TER BLOCK~
15 0 0 90
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
3750 0 0
0
0
10 TER BLOCK~
94 828 493 0 2 5
0 27 44
10 TER BLOCK~
16 0 0 90
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 0 1 0 0 0
0
8778 0 0
0
0
10 TER BLOCK~
94 817 493 0 2 5
0 58 44
10 TER BLOCK~
17 0 0 90
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 0 1 0 0 0
0
538 0 0
0
0
10 TER BLOCK~
94 806 493 0 2 5
0 28 45
10 TER BLOCK~
18 0 0 90
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 0 1 0 0 0
0
6843 0 0
0
0
10 TER BLOCK~
94 795 493 0 2 5
0 59 44
10 TER BLOCK~
19 0 0 90
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 0 1 0 0 0
0
3136 0 0
0
0
10 TER BLOCK~
94 941 493 0 2 5
0 119 50
10 TER BLOCK~
20 0 0 90
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
5950 0 0
0
0
10 TER BLOCK~
94 930 493 0 2 5
0 120 49
10 TER BLOCK~
21 0 0 90
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
5670 0 0
0
0
10 TER BLOCK~
94 919 493 0 2 5
0 121 48
10 TER BLOCK~
22 0 0 90
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
6828 0 0
0
0
10 TER BLOCK~
94 909 493 0 2 5
0 122 47
10 TER BLOCK~
23 0 0 90
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
6735 0 0
0
0
10 TER BLOCK~
94 898 493 0 2 5
0 123 47
10 TER BLOCK~
24 0 0 90
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
8365 0 0
0
0
10 TER BLOCK~
94 887 493 0 2 5
0 124 46
10 TER BLOCK~
25 0 0 90
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
4132 0 0
0
0
10 TER BLOCK~
94 876 493 0 2 5
0 51 32
10 TER BLOCK~
26 0 0 90
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 0 1 0 0 0
0
4551 0 0
0
0
10 TER BLOCK~
94 865 493 0 2 5
0 52 2
10 TER BLOCK~
27 0 0 90
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 0 1 0 0 0
0
3635 0 0
0
0
10 TER BLOCK~
94 854 493 0 2 5
0 25 74
10 TER BLOCK~
28 0 0 90
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 0 1 0 0 0
0
3973 0 0
0
0
10 TER BLOCK~
94 843 493 0 2 5
0 26 50
10 TER BLOCK~
29 0 0 90
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 0 1 0 0 0
0
3851 0 0
0
0
10 TER BLOCK~
94 999 493 0 2 5
0 39 69
10 TER BLOCK~
30 0 0 90
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 0 1 0 0 0
0
8383 0 0
0
0
10 TER BLOCK~
94 988 493 0 2 5
0 40 67
10 TER BLOCK~
31 0 0 90
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 0 1 0 0 0
0
9334 0 0
0
0
10 TER BLOCK~
94 978 493 0 2 5
0 41 68
10 TER BLOCK~
32 0 0 90
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 0 1 0 0 0
0
7471 0 0
0
0
10 TER BLOCK~
94 967 493 0 2 5
0 42 68
10 TER BLOCK~
33 0 0 90
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 0 1 0 0 0
0
3334 0 0
0
0
10 TER BLOCK~
94 956 493 0 2 5
0 43 69
10 TER BLOCK~
34 0 0 90
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 0 1 0 0 0
0
3559 0 0
0
0
10 TER BLOCK~
94 1036 493 0 2 5
0 36 70
10 TER BLOCK~
35 0 0 90
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 0 1 0 0 0
0
984 0 0
0
0
10 TER BLOCK~
94 1025 493 0 2 5
0 37 71
10 TER BLOCK~
36 0 0 90
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 0 1 0 0 0
0
7557 0 0
0
0
10 TER BLOCK~
94 1014 493 0 2 5
0 38 70
10 TER BLOCK~
37 0 0 90
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 0 1 0 0 0
0
3146 0 0
0
0
10 TER BLOCK~
94 1126 493 0 2 5
0 33 60
10 TER BLOCK~
38 0 0 90
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 0 1 0 0 0
0
5687 0 0
0
0
10 TER BLOCK~
94 1115 493 0 2 5
0 34 61
10 TER BLOCK~
39 0 0 90
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 0 1 0 0 0
0
7939 0 0
0
0
10 TER BLOCK~
94 1104 493 0 2 5
0 35 62
10 TER BLOCK~
40 0 0 90
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 0 1 0 0 0
0
3308 0 0
0
0
10 TER BLOCK~
94 1093 493 0 2 5
0 17 63
10 TER BLOCK~
41 0 0 90
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 0 1 0 0 0
0
3408 0 0
0
0
10 TER BLOCK~
94 1082 493 0 2 5
0 18 64
10 TER BLOCK~
42 0 0 90
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 0 1 0 0 0
0
9773 0 0
0
0
10 TER BLOCK~
94 1071 493 0 2 5
0 20 65
10 TER BLOCK~
43 0 0 90
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 0 1 0 0 0
0
691 0 0
0
0
10 TER BLOCK~
94 1061 493 0 2 5
0 24 66
10 TER BLOCK~
44 0 0 90
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 0 1 0 0 0
0
7834 0 0
0
0
10 TER BLOCK~
94 1051 493 0 2 5
0 31 60
10 TER BLOCK~
45 0 0 90
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 0 1 0 0 0
0
3588 0 0
0
0
10 TER BLOCK~
94 1178 243 0 2 5
0 125 4
10 TER BLOCK~
46 0 0 90
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
4528 0 0
0
0
10 TER BLOCK~
94 1188 243 0 2 5
0 126 73
10 TER BLOCK~
47 0 0 90
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
3303 0 0
0
0
10 TER BLOCK~
94 1205 243 0 2 5
0 127 3
10 TER BLOCK~
48 0 0 90
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
9654 0 0
0
0
10 TER BLOCK~
94 1216 243 0 2 5
0 128 72
10 TER BLOCK~
49 0 0 90
0
0
0
0
0
0
0
0
5

0 1 1 1 1 0
0 0 0 512 1 0 0 0
0
9791 0 0
0
0
5 Ter1~
94 856 260 0 1 3
0 67
4 Ter1
50 0 0 90
0
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
4589 0 0
0
0
5 Ter1~
94 866 260 0 1 3
0 48
4 Ter1
51 0 0 90
0
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
964 0 0
0
0
5 Ter1~
94 895 260 0 1 3
0 3
4 Ter1
52 0 0 90
0
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
9151 0 0
0
0
5 Ter1~
94 906 260 0 1 3
0 4
4 Ter1
53 0 0 90
0
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
4745 0 0
0
0
5 Ter1~
94 966 259 0 1 3
0 71
4 Ter1
54 0 0 90
0
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
8433 0 0
0
0
5 Ter1~
94 977 259 0 1 3
0 49
4 Ter1
55 0 0 90
0
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
4221 0 0
0
0
5 Ter1~
94 1001 260 0 1 3
0 72
4 Ter1
56 0 0 90
0
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
8348 0 0
0
0
5 Ter1~
94 1012 260 0 1 3
0 73
4 Ter1
57 0 0 90
0
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
5299 0 0
0
0
5 Ter1~
94 1067 259 0 1 3
0 64
4 Ter1
58 0 0 90
0
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
7393 0 0
0
0
5 Ter1~
94 1077 259 0 1 3
0 50
4 Ter1
59 0 0 90
0
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
6917 0 0
0
0
5 Ter1~
94 1110 259 0 1 3
0 72
4 Ter1
60 0 0 90
0
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
8767 0 0
0
0
5 Ter1~
94 1120 259 0 1 3
0 73
4 Ter1
61 0 0 90
0
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3606 0 0
0
0
5 Ter1~
94 1188 471 0 1 3
0 59
4 Ter1
62 0 0 0
0
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
6970 0 0
0
0
5 Ter1~
94 1188 461 0 1 3
0 52
4 Ter1
63 0 0 0
0
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
343 0 0
0
0
5 Ter1~
94 1188 451 0 1 3
0 8
4 Ter1
64 0 0 0
0
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
7197 0 0
0
0
5 Ter1~
94 1188 441 0 1 3
0 9
4 Ter1
65 0 0 0
0
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3623 0 0
0
0
5 Ter1~
94 1188 431 0 1 3
0 10
4 Ter1
66 0 0 0
0
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
7656 0 0
0
0
5 Ter1~
94 1328 501 0 1 3
0 58
4 Ter1
67 0 0 0
0
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
5365 0 0
0
0
5 Ter1~
94 1328 491 0 1 3
0 51
4 Ter1
68 0 0 0
0
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
4557 0 0
0
0
5 Ter1~
94 1328 481 0 1 3
0 5
4 Ter1
69 0 0 0
0
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3489 0 0
0
0
5 Ter1~
94 1328 471 0 1 3
0 6
4 Ter1
70 0 0 0
0
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
345 0 0
0
0
5 Ter1~
94 1328 461 0 1 3
0 7
4 Ter1
71 0 0 0
0
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3374 0 0
0
0
5 SIP2~
219 191 545 0 2 5
0 43 46
0
0 0 96 180
4 CONN
9 2 37 10
0
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 J
5866 0 0
0
0
11 Contacts:D~
214 331 714 0 10 11
0 77 129 44 0 0 0 0 0 0
1
0
0 0 224 90
6 NORMAL
12 -5 54 3
2 X6
26 -15 40 -7
0
0
18 %D %1 %3 N%D %I %S
0
15 alias:XCONTACTS
4 SIP2
7

0 1 0 2 1 0 2 0
88 0 0 0 1 0 0 0
3 RLY
631 0 0
0
0
11 Contacts:D~
214 357 714 0 10 11
0 77 130 45 0 0 0 0 0 0
1
0
0 0 96 90
6 NORMAL
12 -5 54 3
2 X7
26 -15 40 -7
0
0
18 %D %1 %3 N%D %I %S
0
15 alias:XCONTACTS
4 SIP2
7

0 1 0 2 1 0 2 0
88 0 0 0 1 0 0 0
3 RLY
745 0 0
0
0
5 Ter1~
94 424 511 0 1 3
0 4
4 Ter1
72 0 0 270
0
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
7222 0 0
0
0
5 Ter1~
94 415 511 0 1 3
0 3
4 Ter1
73 0 0 270
0
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
4508 0 0
0
0
5 Ter1~
94 374 512 0 1 3
0 47
4 Ter1
74 0 0 270
0
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3738 0 0
0
0
5 Ter1~
94 364 512 0 1 3
0 77
4 Ter1
75 0 0 270
0
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
91 0 0
0
0
6 CPC14~
94 1823 774 0 14 29
0 16 15 14 13 12 11 131 9 8
7 6 5 132 133
5 CPC14
76 0 4096 90
0
0
0
0
0
0
0
0
29

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 1 2 3 4 5
6 7 8 9 10 11 12 13 14 0
0 0 0 512 1 0 0 0
0
4965 0 0
0
0
6 CPCS9~
94 1819 549 0 1 19
0 0
6 CPCS9~
77 0 4608 90
0
2 U1
-6 -60 8 -52
0
0
0
0
0
0
19

0 1 2 3 4 5 6 7 8 0
1 2 3 4 5 6 7 8 0 0
0 0 0 0 0 0 0 0
0
7791 0 0
0
0
5 CPC9~
94 1826 1077 0 1 19
0 0
5 CPC9~
78 0 4096 0
0
2 U2
75 -4 89 4
0
0
0
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
0 0 0 0 0 0 0 0
1 J
3467 0 0
0
0
5 CPC9~
94 1816 322 0 1 19
0 0
5 CPC9~
79 0 4608 90
0
2 U3
-7 -81 7 -73
0
0
0
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
0 0 0 0 0 0 0 0
0
3907 0 0
0
0
159
5 3 0 0 0 0 0 88 0 0 83 3
1799 322
1799 335
1659 335
2 2 0 0 0 0 0 88 0 0 83 2
1761 322
1659 322
4 2 0 0 0 0 0 88 0 0 82 3
1800 282
1800 270
1680 270
1 1 0 0 0 0 0 88 0 0 82 2
1760 282
1680 282
12 5 0 0 0 0 0 4 6 0 0 7
712 897
757 897
757 712
523 712
523 868
612 868
612 859
9 5 0 0 0 0 0 5 4 0 0 8
692 961
692 951
747 951
747 721
532 721
532 949
612 949
612 937
5 16 0 0 0 0 0 5 4 0 0 8
612 1021
612 1042
541 1042
541 741
737 741
737 934
712 934
712 937
16 10 0 0 0 0 0 4 5 0 0 4
712 937
728 937
728 961
712 961
1 16 0 0 0 0 0 18 6 0 0 8
327 781
321 781
321 833
515 833
515 731
727 731
727 859
712 859
0 8 2 0 0 8320 0 0 0 43 94 3
579 839
548 839
548 561
1 1 3 0 0 4096 0 82 0 0 140 4
415 525
415 533
314 533
314 130
1 1 4 0 0 4096 0 81 0 0 145 4
424 525
424 541
324 541
324 149
1 3 5 0 0 4096 0 75 0 0 19 2
1341 480
1417 480
1 2 6 0 0 4096 0 76 0 0 19 2
1341 470
1417 470
1 1 7 0 0 4096 0 77 0 0 19 2
1341 460
1417 460
12 3 5 0 0 16576 0 85 0 0 19 6
1852 803
1852 791
1881 791
1881 682
1581 682
1581 824
11 2 6 0 0 8384 0 85 0 0 19 4
1826 728
1826 688
1596 688
1596 824
10 1 7 0 0 16576 0 85 0 0 19 6
1825 758
1825 738
1852 738
1852 697
1616 697
1616 824
11 0 1 0 0 4128 0 0 0 0 0 3
1417 450
1417 824
1634 824
1 3 8 0 0 4096 0 70 0 0 25 2
1201 450
1257 450
1 2 9 0 0 4096 0 71 0 0 25 2
1201 440
1257 440
1 1 10 0 0 4224 0 72 0 0 25 2
1201 430
1257 430
9 3 8 0 0 12480 0 85 0 0 25 5
1825 788
1821 788
1821 706
1641 706
1641 847
8 2 9 0 0 12480 0 85 0 0 25 5
1826 818
1816 818
1816 717
1658 717
1658 847
10 0 1 0 0 8224 0 0 0 0 0 3
1257 418
1257 847
1689 847
1 3 11 0 0 4160 0 10 0 0 32 2
1213 1144
1258 1144
1 2 12 0 0 4160 0 11 0 0 32 2
1213 1136
1258 1136
1 1 13 0 0 4160 0 12 0 0 32 2
1213 1126
1258 1126
6 3 11 0 0 8384 0 85 0 0 32 3
1795 758
1695 758
1695 868
5 2 12 0 0 4288 0 85 0 0 32 3
1795 788
1714 788
1714 868
4 1 13 0 0 4288 0 85 0 0 32 3
1796 818
1729 818
1729 868
9 0 1 0 0 8224 0 0 0 0 0 4
1258 1157
1258 868
1738 868
1738 861
1 3 14 0 0 4160 0 15 0 0 39 2
1353 1181
1413 1181
1 2 15 0 0 4160 0 16 0 0 39 2
1353 1171
1413 1171
1 1 16 0 0 4160 0 17 0 0 39 2
1353 1161
1413 1161
3 3 14 0 0 8384 0 85 0 0 39 3
1772 743
1744 743
1744 893
2 2 15 0 0 8384 0 85 0 0 39 3
1772 774
1755 774
1755 893
1 1 16 0 0 8384 0 85 0 0 39 3
1772 803
1768 803
1768 893
8 0 1 0 0 32 0 0 0 0 0 3
1413 1197
1413 893
1779 893
0 0 2 0 0 0 0 0 0 43 42 2
579 859
579 917
1 0 2 0 0 0 0 5 0 0 42 3
591 961
579 961
579 936
3 4 2 0 0 0 0 4 4 0 0 4
591 917
579 917
579 937
591 937
3 4 2 0 0 0 0 6 6 0 0 4
591 839
579 839
579 859
591 859
0 5 17 0 0 8192 0 0 0 51 81 3
611 807
572 807
572 669
0 4 18 0 0 8320 0 0 0 49 81 3
611 886
564 886
564 669
1 5 19 0 0 8320 0 1 5 0 0 4
641 1000
641 1013
612 1013
612 1021
8 2 20 0 0 8192 0 5 1 0 0 4
611 961
611 970
641 970
641 980
5 1 21 0 0 8320 0 4 2 0 0 4
612 937
612 930
641 930
641 917
8 2 18 0 0 0 0 4 2 0 0 4
611 877
611 886
641 886
641 897
5 1 22 0 0 8320 0 6 3 0 0 4
612 859
612 852
641 852
641 841
8 2 17 0 0 0 0 6 3 0 0 4
611 799
611 807
641 807
641 821
0 3 20 0 0 8320 0 0 0 47 81 3
611 970
556 970
556 669
1 1 23 0 0 8320 0 7 18 0 0 3
338 819
327 819
327 781
2 2 24 0 0 4096 0 18 7 0 0 3
367 781
367 819
358 819
1 12 25 0 0 8384 0 14 0 0 96 3
1353 1191
1370 1191
1370 562
1 11 26 0 0 8384 0 9 0 0 96 3
1213 1154
1225 1154
1225 562
1 4 27 0 0 8384 0 13 0 0 112 3
1353 1201
1385 1201
1385 530
1 2 28 0 0 8384 0 8 0 0 112 3
1213 1164
1236 1164
1236 530
0 0 29 0 0 4224 0 0 0 0 0 5
1210 1172
1210 1002
1172 1002
1172 1172
1210 1172
0 0 30 0 0 4224 0 0 0 0 0 5
1349 1209
1349 1032
1312 1032
1312 1209
1349 1209
2 2 24 0 0 8192 0 18 0 0 81 3
367 781
395 781
395 669
1 1 31 0 0 4096 0 19 0 0 81 3
163 741
236 741
236 669
2 7 32 0 0 8320 0 19 0 0 94 5
163 732
179 732
179 610
273 610
273 561
1 8 33 0 0 4224 0 44 0 0 81 2
1124 508
1124 669
1 7 34 0 0 4224 0 45 0 0 81 2
1113 508
1113 669
1 6 35 0 0 4224 0 46 0 0 81 2
1102 508
1102 669
1 5 17 0 0 4224 0 47 0 0 81 2
1091 508
1091 669
1 4 18 0 0 0 0 48 0 0 81 2
1080 508
1080 669
1 3 20 0 0 64 0 49 0 0 81 2
1069 508
1069 669
1 2 24 0 0 4288 0 50 0 0 81 2
1059 508
1059 669
1 1 31 0 0 4288 0 51 0 0 81 2
1049 508
1049 669
1 3 36 0 0 4224 0 41 0 0 82 2
1034 508
1034 622
1 2 37 0 0 4224 0 42 0 0 82 2
1023 508
1023 622
1 1 38 0 0 4224 0 43 0 0 82 2
1012 508
1012 622
1 5 39 0 0 4224 0 36 0 0 83 2
997 508
997 589
1 4 40 0 0 4224 0 37 0 0 83 2
986 508
986 589
1 3 41 0 0 4224 0 38 0 0 83 2
976 508
976 589
1 2 42 0 0 4224 0 39 0 0 83 2
965 508
965 589
1 1 43 0 0 4288 0 40 0 0 83 2
954 508
954 589
1 1 43 0 0 0 0 78 0 0 83 3
195 551
236 551
236 589
7 0 1 0 0 4256 0 0 0 0 0 3
222 669
1698 669
1698 251
6 0 1 0 0 32 0 0 0 0 0 3
785 622
1680 622
1680 266
5 0 1 0 0 32 0 0 0 0 0 3
221 589
1659 589
1659 253
2 3 44 0 0 8320 0 25 79 0 0 6
793 475
793 464
469 464
469 744
331 744
331 732
3 2 45 0 0 12416 0 80 24 0 0 5
357 732
457 732
457 453
804 453
804 475
2 6 46 0 0 4224 0 78 0 0 94 3
195 542
261 542
261 561
1 5 47 0 0 8192 0 83 0 0 94 3
374 526
386 526
386 561
1 4 47 0 0 0 0 83 0 0 94 2
374 526
374 561
1 3 48 0 0 4288 0 57 0 0 95 2
865 245
865 177
1 2 49 0 0 4288 0 61 0 0 95 2
976 244
976 177
1 1 50 0 0 4160 0 65 0 0 95 2
1076 244
1076 177
1 14 51 0 0 8384 0 74 0 0 96 3
1341 490
1360 490
1360 562
1 13 52 0 0 8384 0 69 0 0 96 3
1201 460
1222 460
1222 562
1 0 1 0 0 32 0 0 0 0 0 2
723 561
253 561
1 0 1 0 0 32 0 0 0 0 0 3
725 429
725 177
1091 177
1 0 1 0 0 32 0 0 0 0 0 4
955 429
723 429
723 562
1541 562
1 14 51 0 0 0 0 32 0 0 96 2
874 508
874 562
1 13 52 0 0 0 0 33 0 0 96 2
863 508
863 562
1 12 25 0 0 0 0 34 0 0 96 2
852 508
852 562
1 11 26 0 0 0 0 35 0 0 96 2
841 508
841 562
0 0 53 0 0 4224 0 0 0 0 0 5
1337 508
1337 352
1299 352
1299 508
1337 508
0 0 54 0 0 8320 0 0 0 0 0 5
1196 480
1160 480
1160 322
1196 322
1196 480
0 0 55 0 0 8320 0 0 0 0 0 5
1055 249
1130 249
1130 372
1055 372
1055 249
0 0 56 0 0 8320 0 0 0 0 0 6
957 247
1020 247
1020 337
955 337
955 247
957 247
0 0 57 0 0 8320 0 0 0 0 0 6
845 250
915 250
915 337
846 337
846 250
845 250
1 3 58 0 0 8384 0 73 0 0 112 3
1341 500
1347 500
1347 530
1 4 27 0 0 0 0 22 0 0 112 2
826 508
826 530
1 3 58 0 0 0 0 23 0 0 112 2
815 508
815 530
1 2 28 0 0 0 0 24 0 0 112 2
804 508
804 530
1 1 59 0 0 4096 0 25 0 0 112 2
793 508
793 530
1 1 59 0 0 8384 0 68 0 0 112 3
1201 470
1208 470
1208 530
4 0 1 0 0 32 0 0 0 0 0 2
785 530
1504 530
2 0 44 0 0 0 0 23 0 0 114 2
815 475
815 475
2 2 44 0 0 0 0 25 22 0 0 2
793 475
826 475
2 2 60 0 0 8320 0 51 44 0 0 4
1049 475
1049 469
1124 469
1124 475
2 0 61 0 0 4224 0 45 0 0 0 2
1113 475
1113 469
2 0 62 0 0 4224 0 46 0 0 0 2
1102 475
1102 469
2 0 63 0 0 4224 0 47 0 0 0 2
1091 475
1091 469
2 0 64 0 0 8192 0 48 0 0 122 3
1080 475
1083 475
1083 469
2 0 65 0 0 4224 0 49 0 0 0 2
1069 475
1069 469
2 0 66 0 0 4224 0 50 0 0 0 2
1059 475
1059 469
1 0 64 0 0 16512 0 64 0 0 0 6
1066 244
1066 200
813 200
813 390
1083 390
1083 469
1 0 67 0 0 12416 0 56 0 0 126 6
855 245
855 229
834 229
834 419
986 419
986 469
2 2 50 0 0 4224 0 35 26 0 0 2
841 475
939 475
2 2 68 0 0 8320 0 39 38 0 0 4
965 475
965 469
976 469
976 475
2 0 67 0 0 0 0 37 0 0 0 2
986 475
986 469
2 2 69 0 0 8320 0 36 40 0 0 4
997 475
997 469
954 469
954 475
2 2 70 0 0 8320 0 43 41 0 0 4
1012 475
1012 469
1034 469
1034 475
2 1 71 0 0 8320 0 42 60 0 0 6
1023 475
1023 405
824 405
824 210
965 210
965 244
1 4 72 0 0 4096 0 66 0 0 140 2
1109 244
1109 130
1 4 73 0 0 4096 0 67 0 0 145 2
1119 244
1119 149
1 3 72 0 0 4224 0 62 0 0 140 2
1000 245
1000 130
1 3 73 0 0 4224 0 63 0 0 145 2
1011 245
1011 149
1 2 3 0 0 4096 0 58 0 0 140 2
894 245
894 130
1 2 4 0 0 4096 0 59 0 0 145 2
905 245
905 149
0 4 72 0 0 64 0 0 0 137 140 3
1227 200
1238 200
1238 130
2 3 72 0 0 64 0 55 0 0 140 4
1214 225
1214 220
1227 220
1227 130
0 2 3 0 0 64 0 0 0 139 140 3
1203 209
1215 209
1215 130
2 1 3 0 0 64 0 54 0 0 140 2
1203 225
1203 130
3 0 1 0 0 32 0 0 0 0 0 2
1285 130
289 130
2 4 73 0 0 64 0 53 0 0 145 3
1186 225
1194 225
1194 149
2 1 4 0 0 64 0 52 0 0 145 3
1176 225
1165 225
1165 149
2 3 73 0 0 64 0 53 0 0 145 2
1186 225
1186 149
2 2 4 0 0 64 0 52 0 0 145 2
1176 225
1176 149
2 0 1 0 0 32 0 0 0 0 0 2
1244 149
302 149
2 10 50 0 0 64 0 35 0 0 96 2
841 475
841 429
2 9 74 0 0 4288 0 34 0 0 96 2
852 475
852 429
2 8 2 0 0 64 0 33 0 0 96 2
863 475
863 429
2 7 32 0 0 64 0 32 0 0 96 2
874 475
874 429
2 6 46 0 0 64 0 31 0 0 96 2
885 475
885 429
2 5 47 0 0 4288 0 30 0 0 96 2
896 475
896 429
2 4 47 0 0 64 0 29 0 0 96 2
907 475
907 429
2 3 48 0 0 64 0 28 0 0 96 2
917 475
917 429
2 2 49 0 0 64 0 27 0 0 96 2
928 475
928 429
2 1 50 0 0 64 0 26 0 0 96 2
939 475
939 429
0 0 75 0 0 8320 0 0 0 0 0 6
311 700
311 690
380 690
380 800
311 800
311 700
0 0 76 0 0 8320 0 0 0 0 0 5
350 520
436 520
436 273
350 273
350 520
1 1 77 0 0 16512 0 84 79 0 0 5
364 526
354 526
354 608
331 608
331 696
1 1 77 0 0 0 0 84 80 0 0 4
364 526
364 619
357 619
357 696
20
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
1895 311 1951 335
1899 315 1947 331
6 FEEDER
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 13
1872 535 1984 559
1876 539 1980 555
13 E.STOP SWITCH
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 10
1898 1066 1986 1090
1902 1070 1982 1086
10 AC 110V IN
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 23
1895 768 2087 792
1899 772 2083 788
23 SERVO MOTOR Z1,T1,Z2,T2
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 4
638 955 678 979
642 959 674 975
4 RLY1
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 4
639 870 679 894
643 874 675 890
4 RLY2
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 4
639 792 679 816
643 796 675 812
4 RLY4
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 4
327 750 367 774
331 754 363 770
4 RLY3
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
564 452 596 476
568 456 592 472
3 24V
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
960 408 984 432
964 412 980 428
2 5V
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
992 394 1024 418
996 398 1020 414
3 12V
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
1047 379 1079 403
1051 383 1075 399
3 24V
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
1305 407 1329 431
1309 411 1325 427
2 T2
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
1164 363 1188 387
1168 367 1184 383
2 Z2
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
1178 1050 1202 1074
1182 1054 1198 1070
2 T1
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
1319 1078 1343 1102
1323 1082 1339 1098
2 Z1
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 7
362 384 426 408
366 388 422 404
7 24V/16A
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
858 290 906 314
862 294 902 310
5 5V10A
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
959 287 1015 311
963 291 1011 307
6 12V/5A
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
1066 303 1122 327
1070 307 1118 323
6 24V/5A
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
