CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 280 30 100 9
20 79 780 560
7 5.000 V
7 5.000 V
3 GND
1000 10
24 100 0 1 0
20 Package,Description,
61 C:\PROGRAM FILES\MICROCODE ENGINEERING\CIRCUITMAKER 6\BOM.DAT
0 7
20 79 780 560
145752082 336
1
33 COMMUNICATION
(LASER & FEEDER)

49 MULTITRONIKS
1 FREDERICK ROAD
WARREN, NJ. 07059
10 09-17-1998
0
0
38
5 CON64
94 148 309 0 129 129
0 2 19 64 65 66 67 68 69 70
71 72 73 74 75 76 77 78 79 80
81 82 83 84 85 5 6 86 87 88
7 3 89 90 91 92 31 32 30 29
93 94 22 24 28 27 26 25 23 21
95 53 54 52 51 96 97 43 44 47
48 49 50 46 45 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 -1610612212
5 CON64
1 0 2176 0
0
0
0
0
0
0
0
0
129

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 21 22 23 24 25 26 27 28 29
30 31 32 33 34 35 36 37 38 39
40 41 42 43 44 45 46 47 48 49
50 51 52 53 54 55 56 57 58 59
60 61 62 63 64 1 2 3 4 5
6 7 8 9 10 11 12 13 14 15
16 17 18 19 20 21 22 23 24 25
26 27 28 29 30 31 32 33 34 35
36 37 38 39 40 41 42 43 44 45
46 47 48 49 50 51 52 53 54 55
56 57 58 59 60 61 62 63 64 0
0 0 0 512 1 0 0 0
1 J
8953 0 0
0
0
6 DS8922
94 801 197 0 16 33
0 58 55 19 2 2 2 57 56 43
44 47 48 49 50 46 45
6 DS8922
2 0 2176 0
0
0
0
0
0
0
0
5 DIP16
33

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 1 2 3
4 5 6 7 8 9 10 11 12 13
14 15 16 0
0 0 0 0 1 0 0 0
1 U
4441 0 0
0
0
6 SP232A
94 553 184 0 16 33
0 63 20 62 61 60 59 51 52 57
56 58 55 54 53 2 19
6 SP232A
3 0 4224 0
0
0
0
0
0
0
0
5 DIP16
33

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 1 2 3
4 5 6 7 8 9 10 11 12 13
14 15 16 0
0 0 0 0 1 0 0 0
1 U
3618 0 0
0
0
10 Polar Cap~
219 478 148 0 2 5
0 63 62
0
0 0 832 180
5 0.1uF
-72 -5 -37 3
3 C21
-65 -15 -44 -7
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
6153 0 0
0
0
10 Polar Cap~
219 477 178 0 2 5
0 61 60
0
0 0 832 180
5 0.1uF
-70 -3 -35 5
3 C20
-63 -13 -42 -5
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
5394 0 0
0
0
10 Polar Cap~
219 479 100 0 2 5
0 20 19
0
0 0 832 0
5 0.1uF
-65 -7 -30 1
3 C19
-58 -17 -37 -9
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7734 0 0
0
0
10 Polar Cap~
219 459 234 0 2 5
0 2 59
0
0 0 832 90
5 0.1uF
-53 -6 -18 2
3 C18
-46 -16 -25 -8
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
9914 0 0
0
0
7 Ground~
168 459 268 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3747 0 0
0
0
7 Ground~
168 737 259 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3549 0 0
0
0
7 Ground~
168 892 302 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7931 0 0
0
0
10 Polar Cap~
219 650 119 0 2 5
0 19 2
0
0 0 832 270
5 220uF
-16 -34 19 -26
3 C17
-9 -44 12 -36
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
9325 0 0
0
0
7 Ground~
168 649 138 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8903 0 0
0
0
10 Capacitor~
219 608 232 0 2 5
0 2 19
0
0 0 832 90
6 0.01uF
-48 22 -6 30
3 C16
-37 13 -16 21
0
0
11 %D %1 %2 %V
0
0
6 CAP0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3834 0 0
0
0
7 Ground~
168 608 266 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3363 0 0
0
0
6 DS8922
94 795 471 0 16 33
0 36 33 19 2 2 2 35 34 21
23 25 26 27 28 24 22
6 DS8922
4 0 2176 0
0
0
0
0
0
0
0
5 DIP16
33

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 1 2 3
4 5 6 7 8 9 10 11 12 13
14 15 16 0
0 0 0 0 1 0 0 0
1 U
7668 0 0
0
0
6 SP232A
94 554 458 0 16 33
0 42 38 41 40 39 37 29 30 35
34 36 33 32 31 2 19
6 SP232A
5 0 4224 0
0
0
0
0
0
0
0
5 DIP16
33

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 1 2 3
4 5 6 7 8 9 10 11 12 13
14 15 16 0
0 0 0 0 1 0 0 0
1 U
4718 0 0
0
0
10 Polar Cap~
219 476 422 0 2 5
0 42 41
0
0 0 832 180
5 0.1uF
-79 -5 -44 3
3 C15
-72 -15 -51 -7
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3874 0 0
0
0
10 Polar Cap~
219 474 452 0 2 5
0 40 39
0
0 0 832 180
5 0.1uF
-79 -2 -44 6
3 C14
-72 -12 -51 -4
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
6671 0 0
0
0
10 Polar Cap~
219 452 509 0 2 5
0 2 37
0
0 0 832 90
5 0.1uF
-56 -5 -21 3
3 C13
-49 -15 -28 -7
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3789 0 0
0
0
7 Ground~
168 452 535 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4871 0 0
0
0
7 Ground~
168 741 555 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3750 0 0
0
0
7 Ground~
168 881 571 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8778 0 0
0
0
10 Capacitor~
219 609 515 0 2 5
0 2 19
0
0 0 832 90
6 0.01uF
-49 13 -7 21
3 C12
-33 4 -12 12
0
0
11 %D %1 %2 %V
0
0
6 CAP0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
538 0 0
0
0
7 Ground~
168 609 543 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6843 0 0
0
0
10 Capacitor~
219 707 249 0 2 5
0 2 19
0
0 0 832 90
6 0.01uF
-55 -2 -13 6
3 C11
-45 -12 -24 -4
0
0
11 %D %1 %2 %V
0
0
6 CAP0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3136 0 0
0
0
7 Ground~
168 707 297 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5950 0 0
0
0
10 Polar Cap~
219 491 399 0 2 5
0 38 19
0
0 0 832 0
5 0.1uF
2 -13 37 -5
2 C4
12 -23 26 -15
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
5670 0 0
0
0
10 Capacitor~
219 709 517 0 2 5
0 2 19
0
0 0 832 90
6 0.01uF
-60 -3 -18 5
2 C2
-46 -13 -32 -5
0
0
11 %D %1 %2 %V
0
0
6 CAP0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
6828 0 0
0
0
7 Ground~
168 709 557 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6735 0 0
0
0
7 Ground~
168 64 231 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8365 0 0
0
0
9 Resistor~
219 870 137 0 2 5
0 45 19
0
0 0 864 90
2 1k
-18 -6 -4 2
3 R35
-21 -16 0 -8
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4132 0 0
0
0
9 Resistor~
219 895 139 0 2 5
0 43 19
0
0 0 864 90
2 1k
8 -5 22 3
3 R34
5 -15 26 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4551 0 0
0
0
9 Resistor~
219 869 256 0 3 5
0 2 44 -1
0
0 0 864 90
2 1k
8 -5 22 3
3 R33
5 -15 26 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3635 0 0
0
0
9 Resistor~
219 914 257 0 3 5
0 2 46 -1
0
0 0 864 90
2 1k
8 -5 22 3
3 R32
5 -15 26 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3973 0 0
0
0
9 Resistor~
219 865 407 0 2 5
0 22 19
0
0 0 864 90
2 1k
-21 -5 -7 3
3 R31
-24 -15 -3 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3851 0 0
0
0
9 Resistor~
219 884 406 0 2 5
0 21 19
0
0 0 864 90
2 1k
8 -5 22 3
3 R30
5 -15 26 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8383 0 0
0
0
9 Resistor~
219 863 528 0 3 5
0 2 23 -1
0
0 0 864 90
2 1k
8 -5 22 3
3 R29
5 -15 26 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9334 0 0
0
0
9 Resistor~
219 908 524 0 3 5
0 2 24 -1
0
0 0 864 90
2 1k
8 -5 22 3
3 R28
5 -15 26 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7471 0 0
0
0
87
1 1 2 0 0 0 0 30 1 0 0 3
64 225
64 174
116 174
2 0 19 0 0 4096 0 28 0 0 50 2
709 508
709 456
1 1 2 0 0 0 0 29 28 0 0 2
709 551
709 526
15 0 2 0 0 8320 0 16 0 0 10 4
595 432
625 432
625 531
609 531
2 0 19 0 0 4096 0 23 0 0 50 2
609 506
609 422
0 0 19 0 0 0 0 0 0 87 71 2
626 148
626 100
2 0 19 0 0 0 0 13 0 0 87 2
608 223
608 148
0 2 19 0 0 8320 0 0 1 71 0 5
564 100
564 81
85 81
85 183
116 183
1 2 20 0 0 12416 0 6 3 0 0 4
468 100
453 100
453 158
512 158
1 1 2 0 0 0 0 23 24 0 0 2
609 524
609 537
9 1 21 0 0 8192 0 15 36 0 0 3
827 501
884 501
884 424
0 1 22 0 0 8192 0 0 35 20 0 3
866 438
865 438
865 425
6 0 2 0 0 0 0 15 0 0 37 2
763 483
741 483
15 0 2 0 0 0 0 3 0 0 63 4
594 158
626 158
626 251
608 251
2 0 19 0 0 0 0 25 0 0 87 2
707 240
707 182
1 1 2 0 0 0 0 26 25 0 0 2
707 291
707 258
0 0 19 0 0 0 0 0 0 71 33 2
694 100
694 382
0 49 21 0 0 16512 0 0 1 11 0 5
884 501
884 500
977 500
977 309
180 309
0 48 23 0 0 12416 0 0 1 31 0 4
862 492
969 492
969 318
180 318
16 42 22 0 0 12416 0 15 1 0 0 4
827 438
914 438
914 372
180 372
0 43 24 0 0 12416 0 0 1 30 0 4
908 447
924 447
924 363
180 363
11 47 25 0 0 12416 0 15 1 0 0 4
827 483
961 483
961 327
180 327
12 46 26 0 0 12416 0 15 1 0 0 4
827 474
952 474
952 336
180 336
13 45 27 0 0 12416 0 15 1 0 0 4
827 465
942 465
942 345
180 345
14 44 28 0 0 12416 0 15 1 0 0 4
827 456
933 456
933 354
180 354
7 39 29 0 0 4224 0 16 1 0 0 4
513 482
278 482
278 399
180 399
8 38 30 0 0 4224 0 16 1 0 0 4
513 492
268 492
268 408
180 408
14 36 31 0 0 12416 0 16 1 0 0 6
595 442
647 442
647 565
248 565
248 426
180 426
13 37 32 0 0 12416 0 16 1 0 0 6
595 452
637 452
637 556
258 556
258 417
180 417
15 2 24 0 0 0 0 15 38 0 0 3
827 447
908 447
908 506
10 2 23 0 0 0 0 15 37 0 0 3
827 492
863 492
863 510
2 0 19 0 0 0 0 35 0 0 33 2
865 389
865 382
2 0 19 0 0 0 0 36 0 0 44 4
884 388
884 382
694 382
694 400
1 0 2 0 0 0 0 22 0 0 35 2
881 565
881 553
1 1 2 0 0 0 0 37 38 0 0 4
863 546
863 553
908 553
908 542
5 0 2 0 0 0 0 15 0 0 37 2
763 474
741 474
1 4 2 0 0 0 0 21 15 0 0 3
741 549
741 465
763 465
12 2 33 0 0 4224 0 16 15 0 0 4
595 462
684 462
684 447
763 447
10 8 34 0 0 4224 0 16 15 0 0 4
595 482
725 482
725 501
763 501
9 7 35 0 0 4224 0 16 15 0 0 2
595 492
763 492
11 1 36 0 0 4224 0 16 15 0 0 4
595 472
724 472
724 438
763 438
1 1 2 0 0 0 0 20 19 0 0 2
452 529
452 518
2 6 37 0 0 8320 0 19 16 0 0 3
452 501
452 472
513 472
2 0 19 0 0 0 0 27 0 0 50 4
497 399
497 400
694 400
694 422
2 1 38 0 0 4224 0 16 27 0 0 4
513 432
452 432
452 399
480 399
2 5 39 0 0 12416 0 18 16 0 0 4
464 452
445 452
445 462
513 462
4 1 40 0 0 4224 0 16 18 0 0 2
513 452
481 452
2 3 41 0 0 12416 0 17 16 0 0 4
466 422
444 422
444 442
513 442
1 1 42 0 0 4224 0 16 17 0 0 2
513 422
483 422
16 3 19 0 0 0 0 16 15 0 0 4
595 422
694 422
694 456
763 456
0 57 43 0 0 12416 0 0 1 68 0 6
895 227
983 227
983 18
255 18
255 237
180 237
0 58 44 0 0 12416 0 0 1 67 0 6
868 218
975 218
975 26
245 26
245 228
180 228
0 64 45 0 0 12416 0 0 1 69 0 6
870 164
920 164
920 72
190 72
190 174
180 174
0 63 46 0 0 12416 0 0 1 66 0 6
914 173
930 173
930 64
199 64
199 183
180 183
11 59 47 0 0 12416 0 2 1 0 0 6
833 209
967 209
967 34
237 34
237 219
180 219
12 60 48 0 0 12416 0 2 1 0 0 6
833 200
958 200
958 42
228 42
228 210
180 210
13 61 49 0 0 12416 0 2 1 0 0 6
833 191
948 191
948 49
218 49
218 201
180 201
14 62 50 0 0 12416 0 2 1 0 0 6
833 182
939 182
939 57
208 57
208 192
180 192
7 54 51 0 0 4224 0 3 1 0 0 4
512 208
270 208
270 264
180 264
8 53 52 0 0 4224 0 3 1 0 0 4
512 218
279 218
279 273
180 273
14 51 53 0 0 12416 0 3 1 0 0 4
594 168
645 168
645 291
180 291
13 52 54 0 0 12416 0 3 1 0 0 4
594 178
637 178
637 282
180 282
1 1 2 0 0 0 0 14 13 0 0 2
608 260
608 241
1 2 2 0 0 0 0 12 11 0 0 4
649 132
649 122
649 122
649 126
1 0 19 0 0 0 0 11 0 0 71 2
649 109
649 100
15 2 46 0 0 0 0 2 34 0 0 3
833 173
914 173
914 239
10 2 44 0 0 0 0 2 33 0 0 3
833 218
869 218
869 238
9 1 43 0 0 0 0 2 32 0 0 3
833 227
895 227
895 157
16 1 45 0 0 0 0 2 31 0 0 3
833 164
870 164
870 155
2 0 19 0 0 0 0 31 0 0 71 3
870 119
871 119
871 100
2 2 19 0 0 0 0 32 6 0 0 3
895 121
895 100
485 100
1 0 2 0 0 0 0 10 0 0 73 2
892 296
892 286
1 1 2 0 0 0 0 33 34 0 0 4
869 274
869 286
914 286
914 275
6 0 2 0 0 0 0 2 0 0 76 2
769 209
737 209
5 0 2 0 0 0 0 2 0 0 76 2
769 200
737 200
1 4 2 0 0 0 0 9 2 0 0 3
737 253
737 191
769 191
12 2 55 0 0 12416 0 3 2 0 0 4
594 188
655 188
655 173
769 173
10 8 56 0 0 4224 0 3 2 0 0 4
594 208
719 208
719 227
769 227
9 7 57 0 0 4224 0 3 2 0 0 2
594 218
769 218
11 1 58 0 0 4224 0 3 2 0 0 4
594 198
720 198
720 164
769 164
1 1 2 0 0 0 0 8 7 0 0 2
459 262
459 243
2 6 59 0 0 8320 0 7 3 0 0 3
459 226
459 198
512 198
2 5 60 0 0 12416 0 5 3 0 0 4
467 178
443 178
443 188
512 188
4 1 61 0 0 4224 0 3 5 0 0 2
512 178
484 178
2 3 62 0 0 12416 0 4 3 0 0 4
468 148
443 148
443 168
512 168
1 1 63 0 0 4224 0 3 4 0 0 2
512 148
485 148
16 3 19 0 0 0 0 3 2 0 0 4
594 148
665 148
665 182
769 182
8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
277 559 309 583
281 563 305 579
3 RTS
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
265 539 297 563
269 543 293 559
3 CTS
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
216 384 240 408
220 388 236 404
2 RD
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
269 484 293 508
273 488 289 504
2 TD
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
330 284 362 308
334 288 358 304
3 RTS
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
299 266 331 290
303 270 327 286
3 CTS
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
279 212 303 236
283 216 299 232
2 TD
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
213 247 237 271
217 251 233 267
2 RD
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
