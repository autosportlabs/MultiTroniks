CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
880 1290 30 100 9
0 66 795 572
7 5.000 V
7 5.000 V
3 GND
1000 10
24 100 0 1 0
20 Package,Description,
61 C:\PROGRAM FILES\MICROCODE ENGINEERING\CIRCUITMAKER 6\BOM.DAT
0 7
0 66 795 572
143654930 0
0
0
0
0
0
0
52
5 SIP8~
219 2317 906 0 8 17
0 6 5 4 3 22 21 20 19
0
0 0 608 270
4 CONN
9 2 37 10
4 J14C
-20 13 8 21
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 -1610612604
0 0 0 0 1 0 0 0
1 J
8953 0 0
0
0
5 SIP4~
219 1920 649 0 4 9
0 10 9 8 7
0
0 0 608 692
4 CONN
9 2 37 10
4 J12B
-15 -29 13 -21
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 -1610612604
0 0 0 0 1 0 0 0
1 J
4441 0 0
0
0
5 SIP4~
219 1650 715 0 4 9
0 14 13 12 11
0
0 0 608 90
4 CONN
9 2 37 10
4 J12C
-17 -19 11 -11
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 -1610612604
0 0 0 0 1 0 0 0
1 J
3618 0 0
0
0
5 SIP4~
219 2297 489 0 4 9
0 6 5 4 3
0
0 0 608 512
4 CONN
9 2 37 10
4 J12A
-20 -29 8 -21
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 -1610612604
0 0 0 0 1 0 0 0
1 J
6153 0 0
0
0
5 SIP4~
219 1463 957 0 4 9
0 24 25 26 23
0
0 0 608 270
4 CONN
9 2 37 10
4 J16C
-15 11 13 19
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 -1610612604
0 0 0 0 1 0 0 0
1 J
5394 0 0
0
0
5 SIP4~
219 1437 871 0 4 9
0 22 21 20 19
0
0 0 608 270
4 CONN
9 2 37 10
4 J16A
-18 10 10 18
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 -1610612604
0 0 0 0 1 0 0 0
1 J
7734 0 0
0
0
7 Ground~
168 1930 316 0 1 3
0 2
0
0 0 53344 0
0
4 GND8
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9914 0 0
0
0
5 SIP4~
219 1382 958 0 4 9
0 18 17 16 15
0
0 0 608 270
4 CONN
9 2 37 10
4 J16B
-19 11 9 19
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 -1610612604
0 0 0 0 1 0 0 0
1 J
3747 0 0
0
0
6 CON-64
94 1015 1408 0 129 129
0 2 2 35 94 93 90 92 91 89
88 87 86 85 84 83 82 81 80 79
77 76 75 72 73 74 71 69 70 68
67 67 2 2 66 65 64 63 62 61
60 36 37 38 39 40 41 42 43 44
45 46 47 48 49 50 51 52 53 54
55 56 57 58 59 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 -1610612212
6 CON-64
1 0 4736 0
0
3 J26
-4 -163 17 -155
0
0
0
0
0
6 EURO64
129

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 21 22 23 24 25 26 27 28 29
30 31 32 33 34 35 36 37 38 39
40 41 42 43 44 45 46 47 48 49
50 51 52 53 54 55 56 57 58 59
60 61 62 63 64 1 2 3 4 5
6 7 8 9 10 11 12 13 14 15
16 17 18 19 20 21 22 23 24 25
26 27 28 29 30 31 32 33 34 35
36 37 38 39 40 41 42 43 44 45
46 47 48 49 50 51 52 53 54 55
56 57 58 59 60 61 62 63 64 0
0 0 0 0 1 1 0 0
1 J
3549 0 0
0
0
5 CON20
94 1601 910 0 20 41
0 2 13 11 2 25 23 98 96 2
67 14 12 2 24 26 2 97 95 2
67
5 CON20
2 0 4608 0
0
3 J15
-11 -66 10 -58
0
0
0
0
0
5 IDC20
41

0 1 3 5 7 9 11 13 15 17
19 2 4 6 8 10 12 14 16 18
20 1 3 5 7 9 11 13 15 17
19 2 4 6 8 10 12 14 16 18
20 0
0 0 0 0 1 0 0 0
1 J
7931 0 0
0
0
4 CON4
94 698 219 0 4 9
0 67 35 99 2
4 CON4
3 0 4608 0
4 CON4
-16 -36 12 -28
2 J2
-11 -42 3 -34
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
1 J
9325 0 0
0
0
5 CON20
94 1986 266 0 20 41
0 2 110 2 107 2 104 2 101 2
276 111 109 108 106 105 103 102 100 277
278
5 CON20
4 0 4608 0
0
2 J8
-5 -66 9 -58
0
0
0
0
0
5 IDC20
41

0 1 3 5 7 9 11 13 15 17
19 2 4 6 8 10 12 14 16 18
20 1 3 5 7 9 11 13 15 17
19 2 4 6 8 10 12 14 16 18
20 0
0 0 0 512 1 0 0 0
1 J
8903 0 0
0
0
5 CON10
94 1495 350 0 10 21
0 117 115 114 112 294 2 116 2 113
295
5 CON10
5 0 4608 0
0
2 J5
-19 15 -5 23
0
0
0
0
0
5 IDC10
21

0 2 4 6 8 10 1 3 5 7
9 2 4 6 8 10 1 3 5 7
9 0
0 0 0 512 1 0 0 0
1 A
3834 0 0
0
0
5 CON10
94 2458 933 0 10 21
0 119 120 122 123 296 297 118 298 121
299
5 CON10
6 0 4608 0
0
3 J13
-22 -60 -1 -52
0
0
0
0
0
5 IDC10
21

0 2 4 6 8 10 1 3 5 7
9 2 4 6 8 10 1 3 5 7
9 0
0 0 0 512 1 0 0 0
1 A
3363 0 0
0
0
5 CON10
94 1242 920 0 10 21
0 35 124 65 17 15 2 66 64 18
16
5 CON10
7 0 4608 0
0
3 J17
-20 -61 1 -53
0
0
0
0
0
5 IDC10
21

0 2 4 6 8 10 1 3 5 7
9 2 4 6 8 10 1 3 5 7
9 0
0 0 0 0 1 0 0 0
1 A
7668 0 0
0
0
5 CON50
94 2453 560 0 101 101
0 300 2 6 5 4 3 98 97 301
302 303 304 62 305 306 307 120 308 309
310 119 118 311 312 2 313 2 22 21
20 19 96 95 314 2 315 316 63 317
318 319 123 320 321 322 122 121 323 324
2 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 -1610612324
5 CON50
8 0 2688 0
5 CON50
-18 -132 17 -124
3 J11
-11 -142 10 -134
0
0
0
0
0
5 IDC50
101

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 21 22 23 24 25 26 27 28 29
30 31 32 33 34 35 36 37 38 39
40 41 42 43 44 45 46 47 48 49
50 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 21 22 23 24 25 26 27 28 29
30 31 32 33 34 35 36 37 38 39
40 41 42 43 44 45 46 47 48 49
50 0
0 0 0 512 1 0 0 0
1 J
4718 0 0
0
0
5 DB-37
94 541 1011 0 75 75
0 325 326 127 129 135 132 133 327 328
126 2 329 2 330 2 331 2 332 2
333 334 335 336 337 125 80 90 130 128
134 94 131 86 85 70 83 84 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 -1610612428
5 DB-37
9 0 2560 512
4 DB37
-14 -200 14 -192
3 J18
-17 208 4 216
0
0
0
0
0
6 DB37/M
75

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 21 22 23 24 25 26 27 29 30
31 32 33 34 35 28 37 36 1 2
3 4 5 6 7 8 9 10 11 12
13 14 15 16 17 18 19 20 21 22
23 24 25 26 27 29 30 31 32 33
34 35 28 37 36 0
0 0 0 512 1 0 0 0
1 J
3874 0 0
0
0
5 CON50
94 1155 574 0 101 101
0 375 2 59 58 57 56 376 377 378
379 380 381 71 382 383 384 109 385 386
387 111 110 388 389 2 390 2 55 54
53 52 391 392 393 2 394 395 396 397
398 399 106 400 401 402 108 107 403 404
2 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 -1610612324
5 CON50
10 0 2560 0
5 CON50
-18 -132 17 -124
2 J3
-8 -142 6 -134
0
0
0
0
0
5 IDC50
101

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 21 22 23 24 25 26 27 28 29
30 31 32 33 34 35 36 37 38 39
40 41 42 43 44 45 46 47 48 49
50 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 21 22 23 24 25 26 27 28 29
30 31 32 33 34 35 36 37 38 39
40 41 42 43 44 45 46 47 48 49
50 0
0 0 0 512 1 0 0 0
1 J
6671 0 0
0
0
5 CON50
94 2140 543 0 101 101
0 405 2 51 50 49 48 406 407 408
409 410 411 72 412 413 414 103 415 416
417 105 104 418 419 2 420 2 47 46
45 44 421 422 423 2 424 425 426 427
428 429 100 430 431 432 102 101 433 434
2 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 -1610612324
5 CON50
11 0 2688 0
5 CON50
-18 -132 17 -124
2 J9
-8 -142 6 -134
0
0
0
0
0
5 IDC50
101

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 21 22 23 24 25 26 27 28 29
30 31 32 33 34 35 36 37 38 39
40 41 42 43 44 45 46 47 48 49
50 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 21 22 23 24 25 26 27 28 29
30 31 32 33 34 35 36 37 38 39
40 41 42 43 44 45 46 47 48 49
50 0
0 0 0 512 1 0 0 0
1 J
3789 0 0
0
0
5 DB-37
94 1761 554 0 75 75
0 2 35 435 436 9 7 61 50 48
76 46 44 437 128 126 438 124 67 2
2 35 439 10 8 60 51 49 47 45
440 129 127 441 125 75 2 67 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 -1610612428
5 DB-37
12 0 2688 512
4 DB37
-14 -200 14 -192
2 J7
-7 -210 7 -202
0
0
0
0
0
6 DB37/M
75

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 21 22 23 24 25 26 27 29 30
31 32 33 34 35 28 37 36 1 2
3 4 5 6 7 8 9 10 11 12
13 14 15 16 17 18 19 20 21 22
23 24 25 26 27 29 30 31 32 33
34 35 28 37 36 0
0 0 0 512 1 0 0 0
1 J
4871 0 0
0
0
5 DB-37
94 553 566 0 75 75
0 2 35 99 33 31 29 27 58 56
74 54 52 479 134 132 94 78 67 2
2 35 34 32 30 28 59 57 55 53
480 135 133 131 130 73 2 67 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 -1610612428
5 DB-37
13 0 2688 512
4 DB37
-14 -200 14 -192
2 J1
-8 -201 6 -193
0
0
0
0
0
6 DB37/M
75

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 21 22 23 24 25 26 27 29 30
31 32 33 34 35 28 37 36 1 2
3 4 5 6 7 8 9 10 11 12
13 14 15 16 17 18 19 20 21 22
23 24 25 26 27 29 30 31 32 33
34 35 28 37 36 0
0 0 0 512 1 0 0 0
1 J
3750 0 0
0
0
5 CON50
94 1473 569 0 101 101
0 2 518 30 29 28 27 519 520 521
522 523 524 62 525 526 527 115 528 529
530 117 116 531 532 2 533 2 34 33
32 31 534 535 536 2 537 538 63 539
540 541 112 542 543 544 114 113 545 546
2 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 -1610612488
5 CON50
14 0 2560 0
5 CON50
-18 -132 17 -124
2 J6
-7 -135 7 -127
0
0
0
0
0
5 IDC50
101

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 21 22 23 24 25 26 27 28 29
30 31 32 33 34 35 36 37 38 39
40 41 42 43 44 45 46 47 48 49
50 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 21 22 23 24 25 26 27 28 29
30 31 32 33 34 35 36 37 38 39
40 41 42 43 44 45 46 47 48 49
50 0
0 0 0 512 1 0 0 0
1 J
8778 0 0
0
0
5 SIP8~
219 1246 329 0 8 17
0 55 53 547 548 2 54 52 549
0
0 0 608 90
4 CONN
9 2 37 10
2 J4
-12 -20 2 -12
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 512 1 0 0 0
1 J
538 0 0
0
0
5 SIP8~
219 2239 563 0 8 17
0 47 45 550 551 552 46 44 553
0
0 0 608 90
4 CONN
9 2 37 10
3 J10
-12 -20 9 -12
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 512 1 0 0 0
1 J
6843 0 0
0
0
7 Ground~
168 1816 757 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3136 0 0
0
0
7 Ground~
168 592 765 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5950 0 0
0
0
7 Ground~
168 766 426 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5670 0 0
0
0
7 Ground~
168 723 287 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6828 0 0
0
0
7 Ground~
168 1249 359 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6735 0 0
0
0
7 Ground~
168 1050 647 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8365 0 0
0
0
7 Ground~
168 1310 668 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4132 0 0
0
0
7 Ground~
168 1860 403 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4551 0 0
0
0
7 Ground~
168 2136 701 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3635 0 0
0
0
7 Ground~
168 2415 748 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3973 0 0
0
0
7 Ground~
168 587 1167 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3851 0 0
0
0
7 Ground~
168 909 1294 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8383 0 0
0
0
7 Ground~
168 1436 356 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9334 0 0
0
0
7 Ground~
168 1523 967 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7471 0 0
0
0
7 Ground~
168 1690 965 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3334 0 0
0
0
11 SPDT Relay~
176 834 1290 0 10 11
0 554 555 556 35 93 0 0 0 0
1
0
0 0 4192 512
7 12VSPDT
-25 -35 24 -27
4 RLY1
-14 -45 14 -37
0
0
20 %D %1 %2 %3 %4 %5 %S
0
45 alias:XSPDTRELAY {PULLIN=9.6 RESISTANCE=1000}
4 DIP8
11

0 1 2 3 4 5 1 2 3 4
5 0
88 0 0 512 1 0 0 0
3 RLY
3559 0 0
0
0
5 SIP2~
219 535 1322 0 2 5
0 35 92
0
0 0 608 512
4 CONN
9 2 37 10
3 J19
-16 -20 5 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 J
984 0 0
0
0
5 SIP2~
219 536 1353 0 2 5
0 35 91
0
0 0 608 512
4 CONN
9 2 37 10
3 J20
-17 -20 4 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 J
7557 0 0
0
0
5 SIP4~
219 535 1401 0 4 9
0 89 88 87 67
0
0 0 608 512
4 CONN
9 2 37 10
3 J21
-17 -29 4 -21
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
1 J
3146 0 0
0
0
5 SIP2~
219 535 1456 0 2 5
0 67 82
0
0 0 608 512
4 CONN
9 2 37 10
3 J22
-17 -20 4 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 J
5687 0 0
0
0
5 SIP2~
219 534 1543 0 2 5
0 79 2
0
0 0 608 512
4 CONN
9 2 37 10
3 J24
-17 -20 4 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 J
7939 0 0
0
0
7 Ground~
168 654 1649 0 1 3
0 2
0
0 0 53344 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3308 0 0
0
0
7 Ground~
168 1172 923 0 1 3
0 2
0
0 0 53344 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3408 0 0
0
0
5 SIP3~
219 532 1498 0 3 7
0 67 81 69
0
0 0 608 512
4 CONN
-13 -25 15 -17
3 J23
-14 -25 7 -17
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 J
9773 0 0
0
0
5 SIP4~
219 534 1618 0 4 9
0 78 77 68 2
0
0 0 608 512
4 CONN
9 2 37 10
3 J25
-17 -29 4 -21
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
1 J
691 0 0
0
0
7 Ground~
168 981 1618 0 1 3
0 2
0
0 0 53344 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7834 0 0
0
0
5 SIP8~
219 1326 1448 0 8 17
0 43 42 41 40 39 38 37 36
0
0 0 608 0
4 CONN
9 2 37 10
4 J14A
-14 -47 14 -39
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 0 1 0 0 0
1 J
3588 0 0
0
0
5 SIP8~
219 761 766 0 8 17
0 34 33 32 31 30 29 28 27
0
0 0 608 270
4 CONN
9 2 37 10
4 J14B
35 0 63 8
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 0 1 0 0 0
1 J
4528 0 0
0
0
249
4 0 3 0 0 4224 0 1 0 0 13 2
2319 898
2319 503
0 3 4 0 0 8320 0 0 1 14 0 3
2329 494
2328 494
2328 898
2 0 5 0 0 4224 0 1 0 0 15 2
2337 898
2337 484
0 1 6 0 0 4224 0 0 1 16 0 2
2346 475
2346 898
6 4 7 0 0 8320 0 20 2 0 0 3
1784 636
1784 637
1908 637
24 3 8 0 0 4224 0 20 2 0 0 2
1784 646
1908 646
5 2 9 0 0 8320 0 20 2 0 0 3
1784 656
1784 655
1908 655
23 1 10 0 0 12416 0 20 2 0 0 4
1784 666
1799 666
1799 664
1908 664
3 4 11 0 0 8320 0 10 3 0 0 5
1579 884
1557 884
1557 761
1661 761
1661 724
12 3 12 0 0 8320 0 10 3 0 0 3
1623 874
1652 874
1652 724
2 2 13 0 0 8320 0 10 3 0 0 5
1579 874
1567 874
1567 770
1643 770
1643 724
11 1 14 0 0 8320 0 10 3 0 0 3
1623 864
1634 864
1634 724
4 6 3 0 0 0 0 4 16 0 0 4
2303 503
2406 503
2406 502
2421 502
5 3 4 0 0 0 0 16 4 0 0 4
2421 493
2406 493
2406 494
2303 494
2 4 5 0 0 0 0 4 16 0 0 4
2303 485
2337 485
2337 484
2421 484
3 1 6 0 0 0 0 16 4 0 0 4
2421 475
2346 475
2346 476
2303 476
5 4 15 0 0 4224 0 15 8 0 0 3
1265 920
1366 920
1366 950
10 3 16 0 0 12416 0 15 8 0 0 7
1200 920
1193 920
1193 959
1338 959
1338 930
1375 930
1375 950
4 2 17 0 0 4224 0 15 8 0 0 3
1265 910
1384 910
1384 950
9 1 18 0 0 12416 0 15 8 0 0 7
1200 910
1185 910
1185 969
1348 969
1348 939
1393 939
1393 950
0 8 19 0 0 4096 0 0 1 31 0 2
2283 833
2283 898
7 0 20 0 0 4096 0 1 0 0 37 2
2292 898
2292 823
6 0 21 0 0 4096 0 1 0 0 35 2
2301 898
2301 813
5 0 22 0 0 4096 0 1 0 0 33 2
2310 898
2310 803
1 0 2 0 0 4096 0 7 0 0 28 2
1930 310
1930 300
5 0 2 0 0 4096 0 12 0 0 29 2
1964 260
1930 260
3 0 2 0 0 0 0 12 0 0 29 2
1964 240
1930 240
0 9 2 0 0 0 0 0 12 29 0 3
1930 279
1930 300
1964 300
1 7 2 0 0 8192 0 12 12 0 0 4
1964 220
1930 220
1930 280
1964 280
4 6 23 0 0 8320 0 5 10 0 0 3
1447 949
1447 914
1579 914
4 31 19 0 0 8320 0 6 16 0 0 6
1421 863
1421 833
2549 833
2549 627
2485 627
2485 628
1 14 24 0 0 8320 0 5 10 0 0 5
1474 949
1474 845
1644 845
1644 894
1623 894
1 28 22 0 0 8320 0 6 16 0 0 5
1448 863
1448 803
2516 803
2516 655
2485 655
2 5 25 0 0 8320 0 5 10 0 0 3
1465 949
1465 904
1579 904
2 29 21 0 0 8320 0 6 16 0 0 5
1439 863
1439 813
2528 813
2528 646
2485 646
3 15 26 0 0 16512 0 5 10 0 0 7
1456 949
1456 924
1508 924
1508 993
1643 993
1643 904
1623 904
3 30 20 0 0 8320 0 6 16 0 0 5
1430 863
1430 823
2539 823
2539 637
2485 637
8 0 27 0 0 4096 0 52 0 0 205 2
727 758
727 628
7 0 28 0 0 4096 0 52 0 0 206 2
736 758
736 638
6 0 29 0 0 4096 0 52 0 0 207 2
745 758
745 648
5 0 30 0 0 4096 0 52 0 0 208 2
754 758
754 658
4 0 31 0 0 4096 0 52 0 0 246 2
763 758
763 668
3 0 32 0 0 4096 0 52 0 0 247 2
772 758
772 678
2 0 33 0 0 4096 0 52 0 0 248 2
781 758
781 688
1 0 34 0 0 4096 0 52 0 0 249 2
790 758
790 698
1 0 35 0 0 8192 0 42 0 0 47 3
542 1349
557 1349
557 1318
0 1 35 0 0 4096 0 0 41 118 0 4
884 1248
557 1248
557 1318
541 1318
8 41 36 0 0 4224 0 51 9 0 0 2
1314 1480
1055 1480
42 7 37 0 0 4224 0 9 51 0 0 2
1055 1471
1314 1471
6 43 38 0 0 4224 0 51 9 0 0 2
1314 1462
1055 1462
44 5 39 0 0 4224 0 9 51 0 0 2
1055 1453
1314 1453
4 45 40 0 0 4224 0 51 9 0 0 2
1314 1444
1055 1444
46 3 41 0 0 4224 0 9 51 0 0 2
1055 1435
1314 1435
2 47 42 0 0 4224 0 51 9 0 0 2
1314 1426
1055 1426
48 1 43 0 0 4224 0 9 51 0 0 2
1055 1417
1314 1417
49 0 44 0 0 12416 0 9 0 0 223 5
1055 1408
1226 1408
1226 1274
1985 1274
1985 717
0 50 45 0 0 8320 0 0 9 224 0 5
1995 726
1995 1264
1217 1264
1217 1399
1055 1399
51 0 46 0 0 12416 0 9 0 0 225 5
1055 1390
1208 1390
1208 1255
2004 1255
2004 737
0 52 47 0 0 8320 0 0 9 226 0 5
2011 745
2011 1245
1198 1245
1198 1381
1055 1381
53 0 48 0 0 12416 0 9 0 0 227 5
1055 1372
1189 1372
1189 1236
2020 1236
2020 576
0 54 49 0 0 8320 0 0 9 228 0 5
2028 586
2028 1228
1180 1228
1180 1363
1055 1363
55 0 50 0 0 12416 0 9 0 0 229 5
1055 1354
1172 1354
1172 1219
2067 1219
2067 596
0 56 51 0 0 8320 0 0 9 230 0 5
2057 606
2057 1211
1164 1211
1164 1345
1055 1345
57 0 52 0 0 8320 0 9 0 0 238 5
1055 1336
1141 1336
1141 867
825 867
825 528
0 58 53 0 0 12416 0 0 9 239 0 5
831 538
831 859
1133 859
1133 1327
1055 1327
59 0 54 0 0 8320 0 9 0 0 240 5
1055 1318
1125 1318
1125 850
838 850
838 548
0 60 55 0 0 12416 0 0 9 241 0 5
845 558
845 842
1116 842
1116 1309
1055 1309
61 0 56 0 0 8192 0 9 0 0 242 5
1055 1300
1108 1300
1108 821
852 821
852 588
0 62 57 0 0 12416 0 0 9 243 0 5
859 598
859 814
1100 814
1100 1291
1055 1291
0 63 58 0 0 12416 0 0 9 244 0 5
866 608
866 806
1092 806
1092 1282
1055 1282
0 64 59 0 0 12416 0 0 9 245 0 5
875 618
875 797
1083 797
1083 1273
1055 1273
40 25 60 0 0 12416 0 9 20 0 0 6
1055 1489
1263 1489
1263 1200
1854 1200
1854 626
1784 626
7 39 61 0 0 8320 0 20 9 0 0 6
1784 616
1845 616
1845 1191
1271 1191
1271 1498
1055 1498
0 38 62 0 0 12288 0 0 9 203 0 5
1426 574
1426 760
1287 760
1287 1507
1055 1507
0 37 63 0 0 12288 0 0 9 204 0 5
1532 574
1532 769
1296 769
1296 1516
1055 1516
36 8 64 0 0 8320 0 9 15 0 0 4
1055 1525
1150 1525
1150 901
1200 901
3 35 65 0 0 8320 0 15 9 0 0 4
1265 900
1279 900
1279 1534
1055 1534
7 34 66 0 0 8320 0 15 9 0 0 4
1200 890
1159 890
1159 1543
1055 1543
33 0 2 0 0 12288 0 9 0 0 82 4
1055 1552
1065 1552
1065 1580
981 1580
0 0 67 0 0 12288 0 0 0 101 81 4
594 1489
659 1489
659 1539
971 1539
30 31 67 0 0 0 0 9 9 0 0 4
989 1534
971 1534
971 1543
989 1543
1 32 2 0 0 0 0 50 9 0 0 3
981 1612
981 1552
989 1552
4 0 2 0 0 4096 0 49 0 0 97 2
540 1632
654 1632
3 29 68 0 0 12416 0 49 9 0 0 4
540 1623
762 1623
762 1525
989 1525
3 27 69 0 0 4224 0 48 9 0 0 2
541 1507
989 1507
35 28 70 0 0 8320 0 17 9 0 0 4
564 1023
615 1023
615 1516
989 1516
13 26 71 0 0 8320 0 18 9 0 0 6
1123 579
1066 579
1066 1190
966 1190
966 1498
989 1498
23 13 72 0 0 12416 0 9 19 0 0 6
989 1471
959 1471
959 1180
2094 1180
2094 548
2108 548
24 35 73 0 0 8320 0 9 21 0 0 4
989 1480
687 1480
687 578
576 578
10 25 74 0 0 8320 0 21 9 0 0 4
576 568
696 568
696 1489
989 1489
35 22 75 0 0 12416 0 20 9 0 0 6
1784 566
1836 566
1836 1172
952 1172
952 1462
989 1462
21 10 76 0 0 12416 0 9 20 0 0 6
989 1453
945 1453
945 1162
1827 1162
1827 556
1784 556
1 0 35 0 0 12288 0 15 0 0 118 4
1265 880
1275 880
1275 833
884 833
1 6 2 0 0 0 0 47 15 0 0 3
1172 917
1172 880
1200 880
2 20 77 0 0 12416 0 49 9 0 0 4
540 1614
754 1614
754 1444
989 1444
17 1 78 0 0 8320 0 21 49 0 0 4
576 428
707 428
707 1605
540 1605
1 2 2 0 0 0 0 46 45 0 0 3
654 1643
654 1548
540 1548
1 19 79 0 0 12416 0 45 9 0 0 4
540 1539
650 1539
650 1435
989 1435
18 26 80 0 0 8320 0 9 17 0 0 4
989 1426
677 1426
677 1063
564 1063
2 17 81 0 0 12416 0 48 9 0 0 4
541 1498
641 1498
641 1417
989 1417
1 0 67 0 0 0 0 48 0 0 103 3
541 1489
594 1489
594 1452
2 16 82 0 0 12416 0 44 9 0 0 4
541 1461
633 1461
633 1408
989 1408
1 0 67 0 0 0 0 44 0 0 108 3
541 1452
594 1452
594 1415
15 36 83 0 0 8320 0 9 17 0 0 4
989 1399
666 1399
666 843
564 843
37 14 84 0 0 8320 0 17 9 0 0 4
564 863
656 863
656 1390
989 1390
13 34 85 0 0 8320 0 9 17 0 0 4
989 1381
647 1381
647 883
564 883
33 12 86 0 0 8320 0 17 9 0 0 4
564 903
636 903
636 1372
989 1372
0 4 67 0 0 4096 0 0 43 171 0 3
624 419
624 1415
541 1415
3 11 87 0 0 12416 0 43 9 0 0 4
541 1406
594 1406
594 1363
989 1363
2 10 88 0 0 12416 0 43 9 0 0 4
541 1397
586 1397
586 1354
989 1354
9 1 89 0 0 4224 0 9 43 0 0 4
989 1345
577 1345
577 1388
541 1388
0 3 35 0 0 0 0 0 9 118 0 4
884 1265
939 1265
939 1291
989 1291
27 6 90 0 0 4224 0 17 9 0 0 4
564 1043
932 1043
932 1318
989 1318
8 2 91 0 0 4224 0 9 42 0 0 4
989 1336
569 1336
569 1358
542 1358
2 7 92 0 0 4224 0 41 9 0 0 2
541 1327
989 1327
5 5 93 0 0 4224 0 9 40 0 0 2
989 1309
848 1309
0 4 94 0 0 8192 0 0 9 232 0 4
939 942
976 942
976 1300
989 1300
0 4 35 0 0 4096 0 0 40 170 0 3
884 728
884 1285
848 1285
1 0 2 0 0 0 0 39 0 0 121 2
1690 959
1690 944
16 0 2 0 0 0 0 10 0 0 121 2
1623 914
1690 914
13 19 2 0 0 0 0 10 10 0 0 4
1623 884
1690 884
1690 944
1623 944
1 0 2 0 0 0 0 38 0 0 124 2
1523 961
1523 944
4 0 2 0 0 0 0 10 0 0 124 2
1579 894
1523 894
1 9 2 0 0 0 0 10 10 0 0 4
1579 864
1523 864
1523 944
1579 944
8 0 2 0 0 0 0 13 0 0 126 2
1453 331
1436 331
1 6 2 0 0 0 0 37 13 0 0 3
1436 350
1436 310
1453 310
2 0 2 0 0 0 0 9 0 0 128 2
989 1282
909 1282
1 1 2 0 0 0 0 36 9 0 0 3
909 1288
909 1273
989 1273
0 0 67 0 0 0 0 0 0 130 152 3
1630 955
1716 955
1716 280
10 20 67 0 0 0 0 10 10 0 0 6
1579 954
1575 954
1575 969
1630 969
1630 954
1623 954
33 18 95 0 0 12416 0 16 10 0 0 6
2485 610
2608 610
2608 988
2109 988
2109 934
1623 934
8 32 96 0 0 12416 0 10 16 0 0 6
1579 934
1568 934
1568 976
2597 976
2597 619
2485 619
17 8 97 0 0 12416 0 10 16 0 0 6
1623 924
1666 924
1666 1000
2366 1000
2366 520
2421 520
7 7 98 0 0 12416 0 10 16 0 0 6
1579 924
1534 924
1534 1063
2356 1063
2356 511
2421 511
1 0 2 0 0 4096 0 35 0 0 139 4
587 1161
587 1008
588 1008
588 993
17 0 2 0 0 0 0 17 0 0 139 2
564 873
588 873
15 0 2 0 0 0 0 17 0 0 139 2
564 913
588 913
13 0 2 0 0 0 0 17 0 0 139 2
564 953
588 953
11 19 2 0 0 8192 0 17 17 0 0 4
564 993
588 993
588 833
564 833
1 0 2 0 0 0 0 34 0 0 143 2
2415 742
2415 704
0 50 2 0 0 0 0 0 16 142 0 4
2504 592
2502 592
2502 457
2485 457
0 35 2 0 0 0 0 0 16 143 0 3
2504 665
2504 592
2485 592
0 27 2 0 0 0 0 0 16 144 0 5
2404 672
2404 704
2504 704
2504 664
2485 664
2 25 2 0 0 8192 0 16 16 0 0 4
2421 466
2404 466
2404 673
2421 673
1 0 2 0 0 0 0 33 0 0 148 2
2136 695
2136 682
0 50 2 0 0 0 0 0 19 147 0 3
2188 575
2188 440
2172 440
0 35 2 0 0 0 0 0 19 148 0 3
2188 647
2188 575
2172 575
0 27 2 0 0 0 0 0 19 149 0 5
2086 654
2086 682
2188 682
2188 647
2172 647
2 25 2 0 0 0 0 19 19 0 0 4
2108 449
2086 449
2086 656
2108 656
0 0 35 0 0 12416 0 0 0 151 170 5
1810 707
1809 707
1809 212
884 212
884 213
2 21 35 0 0 0 0 20 20 0 0 4
1784 716
1810 716
1810 706
1784 706
0 0 67 0 0 12416 0 0 0 153 172 4
1828 396
1829 396
1829 280
747 280
37 18 67 0 0 0 0 20 20 0 0 4
1784 406
1828 406
1828 396
1784 396
19 0 2 0 0 0 0 20 0 0 155 3
1784 376
1808 376
1808 386
36 1 2 0 0 0 0 20 32 0 0 3
1784 386
1860 386
1860 397
1 0 2 0 0 0 0 31 0 0 157 3
1310 662
1310 644
1352 644
1 0 2 0 0 8320 0 22 0 0 160 3
1441 466
1352 466
1352 682
50 0 2 0 0 0 0 22 0 0 159 3
1505 466
1521 466
1521 602
0 35 2 0 0 0 0 0 22 160 0 3
1521 674
1521 601
1505 601
25 27 2 0 0 0 0 22 22 0 0 6
1441 682
1352 682
1352 711
1521 711
1521 673
1505 673
1 0 2 0 0 0 0 30 0 0 162 3
1050 641
1050 627
1078 627
2 0 2 0 0 0 0 18 0 0 165 4
1123 480
1078 480
1078 687
1079 687
50 0 2 0 0 0 0 18 0 0 164 3
1187 471
1202 471
1202 607
0 35 2 0 0 0 0 0 18 165 0 3
1202 679
1202 606
1187 606
25 27 2 0 0 0 0 18 18 0 0 6
1123 687
1079 687
1079 711
1202 711
1202 678
1187 678
1 5 2 0 0 0 0 29 23 0 0 3
1249 353
1248 353
1248 338
1 4 2 0 0 0 0 28 11 0 0 3
723 281
723 233
712 233
3 3 99 0 0 8320 0 21 11 0 0 4
576 708
818 708
818 223
712 223
0 21 35 0 0 0 0 0 21 170 0 3
593 729
593 718
576 718
2 2 35 0 0 0 0 11 21 0 0 6
712 213
884 213
884 729
593 729
593 728
576 728
37 0 67 0 0 0 0 21 0 0 172 5
576 418
624 418
624 419
747 419
747 408
18 1 67 0 0 0 0 21 11 0 0 4
576 408
747 408
747 203
712 203
19 0 2 0 0 0 0 21 0 0 174 3
576 388
665 388
665 399
1 36 2 0 0 0 0 27 21 0 0 5
766 420
766 399
665 399
665 398
576 398
1 0 2 0 0 0 0 26 0 0 176 4
592 759
592 755
593 755
593 749
20 1 2 0 0 0 0 21 21 0 0 6
576 738
593 738
593 749
593 749
593 748
576 748
1 0 2 0 0 0 0 25 0 0 178 2
1816 751
1816 735
20 1 2 0 0 0 0 20 20 0 0 4
1784 726
1816 726
1816 736
1784 736
18 42 100 0 0 8320 0 12 19 0 0 4
2008 290
2215 290
2215 512
2172 512
8 47 101 0 0 12416 0 12 19 0 0 6
1964 290
1943 290
1943 342
2205 342
2205 467
2172 467
17 46 102 0 0 8320 0 12 19 0 0 4
2008 280
2196 280
2196 476
2172 476
16 17 103 0 0 8320 0 12 19 0 0 4
2008 270
2077 270
2077 584
2108 584
22 6 104 0 0 8320 0 19 12 0 0 6
2108 629
2038 629
2038 330
1951 330
1951 270
1964 270
15 21 105 0 0 8320 0 12 19 0 0 4
2008 260
2047 260
2047 620
2108 620
14 42 106 0 0 12416 0 12 18 0 0 6
2008 250
2044 250
2044 160
1313 160
1313 543
1187 543
4 47 107 0 0 4224 0 12 18 0 0 4
1964 250
1304 250
1304 498
1187 498
13 46 108 0 0 12416 0 12 18 0 0 6
2008 240
2033 240
2033 170
1295 170
1295 507
1187 507
17 12 109 0 0 12416 0 18 12 0 0 6
1123 615
1086 615
1086 182
2023 182
2023 230
2008 230
2 22 110 0 0 4224 0 12 18 0 0 4
1964 230
1095 230
1095 660
1123 660
21 11 111 0 0 12416 0 18 12 0 0 6
1123 651
1105 651
1105 191
2014 191
2014 220
2008 220
4 42 112 0 0 8320 0 13 22 0 0 4
1518 340
1559 340
1559 538
1505 538
9 47 113 0 0 12416 0 13 22 0 0 6
1453 340
1416 340
1416 397
1541 397
1541 493
1505 493
3 46 114 0 0 8320 0 13 22 0 0 4
1518 330
1550 330
1550 502
1505 502
2 17 115 0 0 16512 0 13 22 0 0 6
1518 320
1530 320
1530 369
1362 369
1362 610
1441 610
7 22 116 0 0 8320 0 13 22 0 0 4
1453 320
1371 320
1371 655
1441 655
1 21 117 0 0 16512 0 13 22 0 0 6
1518 310
1540 310
1540 379
1380 379
1380 646
1441 646
22 7 118 0 0 8320 0 16 14 0 0 4
2421 646
2374 646
2374 903
2416 903
21 1 119 0 0 8320 0 16 14 0 0 6
2421 637
2384 637
2384 872
2483 872
2483 893
2481 893
17 2 120 0 0 8320 0 16 14 0 0 6
2421 601
2394 601
2394 864
2494 864
2494 903
2481 903
47 9 121 0 0 8320 0 16 14 0 0 6
2485 484
2588 484
2588 854
2404 854
2404 923
2416 923
46 3 122 0 0 8320 0 16 14 0 0 4
2485 493
2578 493
2578 913
2481 913
42 4 123 0 0 8320 0 16 14 0 0 4
2485 529
2568 529
2568 923
2481 923
13 13 62 0 0 20608 0 22 16 0 0 8
1441 574
1425 574
1425 388
1618 388
1618 353
2381 353
2381 565
2421 565
38 38 63 0 0 12416 0 16 22 0 0 6
2485 565
2559 565
2559 846
1726 846
1726 574
1505 574
7 6 27 0 0 4224 0 21 22 0 0 6
576 628
996 628
996 378
1323 378
1323 511
1441 511
25 5 28 0 0 4224 0 21 22 0 0 6
576 638
1004 638
1004 388
1400 388
1400 502
1441 502
6 4 29 0 0 4224 0 21 22 0 0 6
576 648
1013 648
1013 398
1409 398
1409 493
1441 493
24 3 30 0 0 4224 0 21 22 0 0 6
576 658
1022 658
1022 407
1418 407
1418 484
1441 484
7 0 44 0 0 0 0 24 0 0 223 2
2259 572
2259 611
6 0 46 0 0 0 0 24 0 0 225 3
2250 572
2249 572
2249 629
2 0 45 0 0 0 0 24 0 0 224 2
2214 572
2214 620
1 0 47 0 0 0 0 24 0 0 226 3
2205 572
2204 572
2204 638
0 7 52 0 0 0 0 0 23 238 0 3
1245 642
1266 642
1266 338
0 6 54 0 0 0 0 0 23 240 0 3
1225 661
1257 661
1257 338
0 2 53 0 0 0 0 0 23 239 0 2
1221 651
1221 338
0 1 55 0 0 0 0 0 23 241 0 2
1212 669
1212 338
2 17 124 0 0 12416 0 15 20 0 0 6
1265 890
1304 890
1304 779
1948 779
1948 416
1784 416
34 25 125 0 0 12416 0 20 17 0 0 4
1784 426
1865 426
1865 1083
564 1083
15 10 126 0 0 12416 0 20 17 0 0 4
1784 456
1874 456
1874 1013
564 1013
32 3 127 0 0 12416 0 20 17 0 0 4
1784 466
1958 466
1958 1153
564 1153
14 29 128 0 0 12416 0 20 17 0 0 5
1784 476
1968 476
1968 984
564 984
564 983
31 4 129 0 0 12416 0 20 17 0 0 4
1784 486
1976 486
1976 1133
564 1133
12 31 44 0 0 0 0 20 19 0 0 6
1784 516
1985 516
1985 717
2259 717
2259 611
2172 611
29 30 45 0 0 0 0 20 19 0 0 6
1784 526
1995 526
1995 727
2214 727
2214 620
2172 620
11 29 46 0 0 0 0 20 19 0 0 6
1784 536
2004 536
2004 737
2249 737
2249 629
2172 629
28 28 47 0 0 0 0 20 19 0 0 6
1784 546
2011 546
2011 745
2204 745
2204 638
2172 638
9 6 48 0 0 0 0 20 19 0 0 4
1784 576
2020 576
2020 485
2108 485
27 5 49 0 0 0 0 20 19 0 0 4
1784 586
2029 586
2029 476
2108 476
8 4 50 0 0 0 0 20 19 0 0 4
1784 596
2067 596
2067 467
2108 467
26 3 51 0 0 0 0 20 19 0 0 4
1784 606
2057 606
2057 458
2108 458
34 28 130 0 0 8320 0 21 17 0 0 4
576 438
949 438
949 1003
564 1003
16 31 94 0 0 8320 0 21 17 0 0 4
576 448
939 448
939 943
564 943
33 32 131 0 0 8320 0 21 17 0 0 4
576 458
930 458
930 923
564 923
6 15 132 0 0 8320 0 17 21 0 0 4
564 1093
920 1093
920 468
576 468
32 7 133 0 0 8320 0 21 17 0 0 4
576 478
910 478
910 1073
564 1073
30 14 134 0 0 8320 0 17 21 0 0 4
564 963
903 963
903 488
576 488
31 5 135 0 0 8320 0 21 17 0 0 4
576 498
893 498
893 1113
564 1113
12 31 52 0 0 0 0 21 18 0 0 6
576 528
957 528
957 779
1245 779
1245 642
1187 642
29 30 53 0 0 0 0 21 18 0 0 6
576 538
967 538
967 769
1234 769
1234 651
1187 651
11 29 54 0 0 0 0 21 18 0 0 6
576 548
977 548
977 761
1225 761
1225 660
1187 660
28 28 55 0 0 0 0 21 18 0 0 6
576 558
986 558
986 752
1212 752
1212 669
1187 669
9 6 56 0 0 4224 0 21 18 0 0 4
576 588
1057 588
1057 516
1123 516
27 5 57 0 0 0 0 21 18 0 0 4
576 598
1048 598
1048 507
1123 507
8 4 58 0 0 0 0 21 18 0 0 4
576 608
1039 608
1039 498
1123 498
26 3 59 0 0 0 0 21 18 0 0 4
576 618
1030 618
1030 489
1123 489
5 31 31 0 0 12416 0 21 22 0 0 6
576 668
1017 668
1017 743
1570 743
1570 637
1505 637
23 30 32 0 0 12416 0 21 22 0 0 6
576 678
1027 678
1027 732
1560 732
1560 646
1505 646
4 29 33 0 0 12416 0 21 22 0 0 6
576 688
1037 688
1037 721
1551 721
1551 655
1505 655
22 28 34 0 0 12416 0 21 22 0 0 6
576 698
1009 698
1009 789
1542 789
1542 664
1505 664
21
-15 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 8
404 1530 485 1555
408 1534 480 1551
8 RESET SW
-15 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 9
401 1595 491 1620
405 1599 486 1616
9 E.STOP SW
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
1185 835 1281 859
1189 839 1277 855
11 Y INTERFACE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
2408 394 2488 418
2412 398 2484 414
9 XY ROTARY
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
2076 397 2116 421
2080 401 2112 417
4 Z2T2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1448 412 1504 436
1452 416 1500 432
6 XY LIN
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1130 407 1170 431
1134 411 1166 427
4 Z1T1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
2190 521 2278 545
2194 525 2274 541
10 LASER ENC2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
1201 276 1289 300
1205 280 1285 296
10 LASER ENC1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
1473 841 1585 865
1477 845 1581 861
13 AC MOTOR ENC.
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 19
2379 940 2539 964
2383 944 2535 960
19  MOTOR DRIVE RORARY
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 15
1428 276 1556 300
1432 280 1552 296
15 MOTOR DRIVE LIN
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
469 1224 573 1248
473 1228 569 1244
12 TO DIO BOARD
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
440 1311 512 1335
444 1315 508 1331
8 DOOR SW1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
437 1340 509 1364
441 1344 505 1360
8 DOOR SW2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
410 1384 506 1408
414 1388 502 1404
11 TOWER LIGHT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
399 1440 503 1464
403 1444 499 1460
12 X,Y SERVO ON
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
401 1478 497 1522
405 1482 493 1514
21 Z1,T1,Z2,T2
SERO ON
-15 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 17
1818 188 1980 213
1822 192 1975 209
17 Z1,T1,Z2,T2 DRIVE
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 11
1609 676 1693 696
1613 680 1690 694
11 AC X ROTARY
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 8
1885 668 1948 688
1889 672 1945 686
8 X ROTARY
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
