CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 40 9
20 78 780 559
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
65 C:\PROGRAM FILES\MICROCODE ENGINEERING\CIRCUITMAKER 6 PRO\BOM.DAT
0 7
20 78 780 559
146341906 0
0
6 Title:
5 Name:
10 10-15-1998
0
4 LVX2
4
2 SC
94 724 369 0 1 3
0 0
2 SC
9 0 0 0
0
2 U4
-10 -45 4 -37
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 0 0 0 0
1 J
8953 0 0
0
0
2 SC
94 666 370 0 1 3
0 0
2 SC
8 0 0 0
0
2 U3
-10 -45 4 -37
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 0 0 0 0
1 J
4441 0 0
0
0
6 CIRCLE
94 384 240 0 1 3
0 0
6 CIRCLE
7 0 0 0
0
2 U2
-14 -63 0 -55
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
1 J
3618 0 0
0
0
6 CIRCLE
94 277 238 0 1 3
0 0
6 CIRCLE
6 0 0 0
0
2 U1
-14 -63 0 -55
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
1 J
6153 0 0
0
0
35
0 0 0 0 0 0 0 0 0 0 0 2
794 248
822 248
0 0 0 0 0 0 0 0 0 0 0 2
796 212
824 212
0 0 0 0 0 0 0 0 0 0 0 5
55 483
481 483
481 576
55 576
55 477
0 0 0 0 0 0 0 0 0 0 0 4
563 304
563 599
454 599
454 576
0 0 0 0 0 0 0 0 0 0 0 4
426 459
426 441
447 441
447 460
0 0 0 0 0 0 0 0 0 0 0 4
741 459
741 441
762 441
762 460
0 0 0 0 0 0 0 0 0 0 0 4
173 459
173 441
194 441
194 460
0 0 0 0 0 0 0 0 0 0 0 4
89 461
89 468
833 468
833 461
0 0 0 0 0 0 0 0 0 0 0 5
799 412
821 412
821 436
799 436
799 412
0 0 0 0 0 0 0 0 0 0 0 6
799 344
821 344
821 367
798 367
798 344
799 344
0 0 0 0 0 0 0 0 0 0 0 5
795 177
823 177
823 287
795 287
795 177
0 0 2 0 0 0 0 0 0 0 0 5
624 308
663 308
663 321
624 321
624 308
0 0 3 0 0 0 0 0 0 0 0 6
554 273
521 273
521 261
556 261
556 273
554 273
0 0 4 0 0 0 0 0 0 0 0 6
565 278
551 278
551 304
605 304
605 278
565 278
0 0 5 0 0 0 0 0 0 0 0 5
594 286
599 286
599 292
594 292
594 286
0 0 6 0 0 0 0 0 0 0 0 5
575 286
581 286
581 292
575 292
575 286
0 0 7 0 0 0 0 0 0 0 0 5
558 286
563 286
563 292
558 292
558 286
0 0 8 0 0 0 0 0 0 0 0 2
551 298
606 298
0 0 9 0 0 0 0 0 0 0 0 5
659 286
664 286
664 292
659 292
659 286
0 0 10 0 0 0 0 0 0 0 0 5
640 286
646 286
646 292
640 292
640 286
0 0 11 0 0 0 0 0 0 0 0 5
623 286
628 286
628 292
623 292
623 286
0 0 12 0 0 0 0 0 0 0 0 2
616 298
671 298
0 0 13 0 0 0 0 0 0 0 0 6
624 278
671 278
671 303
616 303
616 278
624 278
0 0 14 0 0 0 0 0 0 0 0 4
654 184
675 184
675 250
654 250
0 0 15 0 0 0 0 0 0 0 0 4
624 183
604 183
604 250
624 250
0 0 16 0 0 0 0 0 0 0 0 5
624 171
654 171
654 264
624 264
624 171
0 0 17 0 0 0 0 0 0 0 0 2
250 418
330 418
0 0 18 0 0 0 0 0 0 0 0 2
250 356
330 356
0 0 19 0 0 0 0 0 0 0 0 6
331 423
331 348
250 348
250 425
331 425
331 423
0 0 20 0 0 0 0 0 0 0 0 2
380 419
459 419
0 0 21 0 0 0 0 0 0 0 0 2
379 356
459 356
0 0 22 0 0 0 0 0 0 0 0 5
380 348
380 426
459 426
459 348
380 348
0 0 23 0 0 0 0 0 0 0 0 5
366 336
474 336
474 441
366 441
366 336
0 0 24 0 0 0 0 0 0 0 0 5
231 334
349 334
349 441
231 441
231 334
0 0 25 0 0 0 0 0 0 0 0 5
89 155
832 155
832 461
89 461
89 155
20
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
624 302 662 325
629 307 659 322
4 230V
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
520 254 558 277
525 259 555 274
4 115V
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
316 222 332 245
321 227 329 242
1 +
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
207 221 223 244
212 226 220 241
1 +
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
654 384 670 407
659 389 667 404
1 +
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
713 383 729 406
718 388 726 403
1 +
-19 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 93
63 504 479 591
68 509 473 572
93 PLEASE UNPLUG THE WIRES FROM THIS
CONNECTOR AND PLUG IT TO THE HEADER
WHICH IS LABELED 230V
-16 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 14
253 363 323 418
259 368 319 408
14 TRANSF
ORMER
-16 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 14
385 359 455 414
391 364 451 404
14 TRANSF
ORMER
-16 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 14
605 191 675 246
611 196 671 236
14 TRANSF
ORMER
-16 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 10
266 281 376 311
272 284 372 304
10 CAPACITORS
-16 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 10
638 400 748 430
644 403 744 423
10 CAPACITORS
-16 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
798 180 818 210
805 185 815 205
1 G
-16 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
799 217 819 247
805 222 815 242
1 L
-16 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
799 253 819 283
805 258 815 278
1 N
-16 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 4
819 409 869 439
825 414 865 434
4 +OUT
-16 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 4
819 340 869 370
825 345 865 365
4 -OUT
-16 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 9
830 375 930 405
836 380 926 400
9 24VDC/16A
-16 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
830 219 890 249
836 224 886 244
5 AC IN
-16 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 27
108 484 388 514
115 489 385 509
27 IN THE CASE OF 230VAC INPUT
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
